* NGSPICE file created from top_3d_jscan.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt top_3d_jscan VGND VPWR fault_flag reset_n scan_clk scan_in test_enable
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_294_ GTC.mode_sel\[0\] VGND VGND VPWR VPWR _294_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ clknet_2_3__leaf_scan_clk _037_ net10 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_200_ _097_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
X_131_ _054_ _055_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout7 net1 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 TIER1.MSS.scan_chain\[1\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 TIER1.MSS.scan_chain\[6\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold52 GTC.shift_en VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ GTC.col_addr\[3\] VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_276_ clknet_2_0__leaf_scan_clk _036_ VGND VGND VPWR VPWR TIER2.PRAS.scan_out sky130_fd_sc_hd__dfxtp_1
X_130_ _049_ GTC.cluster_sel\[0\] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nand2_1
X_259_ clknet_2_3__leaf_scan_clk _019_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8 net10 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
Xhold42 TIER2.MSS.scan_chain\[4\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _080_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 _113_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ GTC.col_addr\[2\] VGND VGND VPWR VPWR _292_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_275_ clknet_2_3__leaf_scan_clk _035_ net9 VGND VGND VPWR VPWR TIER3.LC.scan_out
+ sky130_fd_sc_hd__dfrtp_1
X_258_ clknet_2_3__leaf_scan_clk _018_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_189_ net2 net37 _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout9 net10 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
Xhold43 TIER2.MSS.scan_chain\[1\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 TIER2.MSS.scan_chain\[2\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold10 GTC.col_addr\[0\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 GTC.tier_sel\[2\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ GTC.col_addr\[1\] VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__buf_2
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_274_ clknet_2_0__leaf_scan_clk _034_ net6 VGND VGND VPWR VPWR GTC.misr_t2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_257_ clknet_2_3__leaf_scan_clk _017_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_188_ _051_ _062_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__nand2_4
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold22 TIER1.MSS.scan_chain\[5\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _095_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 TIER2.LC.scan_out VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 GTC.tier_sel\[0\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_290_ TIER1.tier_sel\[0\] VGND VGND VPWR VPWR _290_/X sky130_fd_sc_hd__buf_2
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_273_ clknet_2_1__leaf_scan_clk _033_ net7 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_256_ clknet_2_3__leaf_scan_clk _016_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_187_ _090_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
X_239_ _050_ net21 _102_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__a21bo_1
Xhold34 TIER1.MSS.scan_chain\[2\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 TIER2.MSS.scan_chain\[3\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 _079_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 GTC.col_addr\[1\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ clknet_2_1__leaf_scan_clk _032_ net6 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_255_ clknet_2_3__leaf_scan_clk _015_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_186_ net28 _084_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_169_ _078_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
X_238_ _050_ net18 _052_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold24 TIER1.MSS.scan_chain\[4\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 _076_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 TIER3.MSS.scan_chain\[5\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 TIER3.PRAS.scan_out VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_271_ clknet_2_1__leaf_scan_clk _031_ net6 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_254_ clknet_2_1__leaf_scan_clk _014_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_185_ net8 _052_ _066_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_168_ net34 net32 _072_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_237_ _050_ net31 _051_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21o_1
Xhold25 TIER2.MSS.scan_chain\[5\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 TIER1.LC.scan_out VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 TIER3.MSS.scan_chain\[2\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold14 TIER2.PRAS.scan_out VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ clknet_2_1__leaf_scan_clk _030_ net6 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ _088_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
X_253_ clknet_2_1__leaf_scan_clk _013_ net6 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_167_ _077_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__clkbuf_1
X_236_ net14 _119_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold37 TIER3.MSS.scan_chain\[0\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _098_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 GTC.col_addr\[2\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 TIER3.MSS.scan_chain\[4\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
X_219_ net47 net48 _108_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__mux2_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_252_ clknet_2_1__leaf_scan_clk _012_ net9 VGND VGND VPWR VPWR TIER1.LC.scan_out
+ sky130_fd_sc_hd__dfrtp_1
X_183_ net54 net2 _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ _065_ TIER3.LC.scan_out _117_ _118_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o211a_1
X_166_ net59 net34 _072_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold16 TIER1.MSS.scan_chain\[0\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 TIER1.MSS.scan_chain\[3\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 TIER2.MSS.scan_chain\[0\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 TIER3.MSS.scan_chain\[1\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _109_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__clkbuf_1
X_149_ _066_ GTC.mode_sel\[1\] _063_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ GTC.mode_sel\[0\] _051_ GTC.mode_sel\[1\] VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__and3b_1
X_251_ clknet_2_2__leaf_scan_clk net19 net8 VGND VGND VPWR VPWR TIER1.tier_sel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_165_ net45 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_234_ TIER3.MSS.scan_chain\[7\] _061_ _081_ TIER3.PRAS.scan_out VGND VGND VPWR VPWR
+ _118_ sky130_fd_sc_hd__o22a_1
Xhold17 _074_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 TIER2.MSS.scan_chain\[6\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 TIER3.MSS.scan_chain\[6\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
X_217_ net2 net47 _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_148_ _065_ GTC.mode_sel\[0\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__and2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ clknet_2_2__leaf_scan_clk _000_ net8 VGND VGND VPWR VPWR TIER1.tier_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_181_ _086_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_302_ net2 VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__buf_2
X_164_ net44 TIER1.MSS.scan_chain\[3\] _072_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_233_ _049_ GTC.tier_sel\[2\] GTC.capture_en VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__and3_1
Xhold18 TIER1.PRAS.scan_out VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _116_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_147_ GTC.mode_sel\[1\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__inv_2
X_216_ _107_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__buf_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout10 net1 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
X_180_ net23 _084_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_163_ _075_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__clkbuf_1
X_301_ net3 VGND VGND VPWR VPWR _301_/X sky130_fd_sc_hd__buf_2
XFILLER_0_5_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_232_ net39 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold19 TIER3.MSS.scan_chain\[3\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_215_ _061_ _102_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__or2_1
X_146_ _064_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_129_ _049_ GTC.cluster_sel\[0\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_162_ net51 net44 _072_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_300_ GTC.shift_en VGND VGND VPWR VPWR _300_/X sky130_fd_sc_hd__buf_2
X_231_ net38 TIER3.MSS.scan_chain\[7\] _108_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__mux2_1
Xinput1 reset_n VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _106_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__clkbuf_1
X_145_ _062_ GTC.mode_sel\[0\] _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _049_ net16 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_scan_clk clknet_0_scan_clk VGND VGND VPWR VPWR clknet_2_3__leaf_scan_clk
+ sky130_fd_sc_hd__clkbuf_16
X_161_ net27 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__clkbuf_1
X_230_ _115_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__clkbuf_1
Xinput2 scan_in VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_144_ GTC.col_addr\[3\] _059_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__nand2_1
X_213_ net24 _084_ _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_127_ _053_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2__f_scan_clk clknet_0_scan_clk VGND VGND VPWR VPWR clknet_2_2__leaf_scan_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_160_ net26 TIER1.MSS.scan_chain\[1\] _072_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_289_ GTC.col_addr\[0\] VGND VGND VPWR VPWR _289_/X sky130_fd_sc_hd__buf_2
Xinput3 test_enable VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ net5 _051_ _066_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__and3_1
X_143_ _061_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_126_ GTC.capture_en net62 _049_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1__f_scan_clk clknet_0_scan_clk VGND VGND VPWR VPWR clknet_2_1__leaf_scan_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ clknet_2_2__leaf_scan_clk _048_ net8 VGND VGND VPWR VPWR GTC.tier_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _104_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
X_142_ GTC.mode_sel\[1\] GTC.mode_sel\[0\] VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_scan_clk clknet_0_scan_clk VGND VGND VPWR VPWR clknet_2_0__leaf_scan_clk
+ sky130_fd_sc_hd__clkbuf_16
X_125_ _050_ GTC.tier_sel\[2\] net18 _052_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_287_ clknet_2_2__leaf_scan_clk _047_ net8 VGND VGND VPWR VPWR GTC.tier_sel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ net17 _059_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__xor2_1
X_210_ net2 net60 _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_124_ net3 GTC.tier_sel\[0\] VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__and2_2
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_286_ clknet_2_2__leaf_scan_clk _046_ net8 VGND VGND VPWR VPWR GTC.tier_sel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ _059_ _060_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nor2_1
X_269_ clknet_2_1__leaf_scan_clk _029_ net6 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_123_ _050_ GTC.tier_sel\[0\] _051_ net31 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_285_ clknet_2_0__leaf_scan_clk net15 net5 VGND VGND VPWR VPWR GTC.misr_t3 sky130_fd_sc_hd__dfrtp_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_268_ clknet_2_1__leaf_scan_clk _028_ net7 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_199_ net52 net35 _091_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_122_ net3 GTC.tier_sel\[1\] VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__and2_2
XFILLER_0_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ clknet_2_2__leaf_scan_clk _044_ net10 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ clknet_2_1__leaf_scan_clk _027_ net7 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_198_ _096_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_121_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ clknet_2_2__leaf_scan_clk _043_ net8 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ net55 net52 _091_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__mux2_1
X_266_ clknet_2_1__leaf_scan_clk _026_ net6 VGND VGND VPWR VPWR TIER2.MSS.scan_chain\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_120_ net3 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_249_ clknet_2_0__leaf_scan_clk _011_ net7 VGND VGND VPWR VPWR GTC.mode_sel\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 GTC.misr_t2 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_scan_clk scan_clk VGND VGND VPWR VPWR clknet_0_scan_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ clknet_2_2__leaf_scan_clk _042_ net8 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ net43 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
X_265_ clknet_2_2__leaf_scan_clk _025_ VGND VGND VPWR VPWR TIER1.PRAS.scan_out sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ _049_ GTC.tier_sel\[2\] net8 _066_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__and4_1
X_248_ clknet_2_0__leaf_scan_clk _010_ net6 VGND VGND VPWR VPWR GTC.mode_sel\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 GTC.misr_t1 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_281_ clknet_2_2__leaf_scan_clk _041_ net8 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ net42 TIER2.MSS.scan_chain\[3\] _091_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__mux2_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ clknet_2_1__leaf_scan_clk _024_ net6 VGND VGND VPWR VPWR TIER2.LC.scan_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_247_ clknet_2_0__leaf_scan_clk _009_ net5 VGND VGND VPWR VPWR GTC.col_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_178_ GTC.col_addr\[0\] GTC.col_addr\[2\] VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 GTC.cluster_sel\[1\] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_280_ clknet_2_3__leaf_scan_clk _040_ net10 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ _094_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ clknet_2_2__leaf_scan_clk _023_ VGND VGND VPWR VPWR TIER3.PRAS.scan_out sky130_fd_sc_hd__dfxtp_1
X_246_ clknet_2_0__leaf_scan_clk _008_ net5 VGND VGND VPWR VPWR GTC.col_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_177_ net12 _083_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__xor2_1
X_229_ net56 net38 _108_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 GTC.misr_t3 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ net53 net42 _091_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__mux2_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ clknet_2_1__leaf_scan_clk _022_ net6 VGND VGND VPWR VPWR GTC.misr_t1 sky130_fd_sc_hd__dfrtp_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_245_ clknet_2_0__leaf_scan_clk _007_ net5 VGND VGND VPWR VPWR GTC.col_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_176_ _065_ TIER1.LC.scan_out _052_ _082_ GTC.capture_en VGND VGND VPWR VPWR _083_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ _073_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
X_228_ _114_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 _045_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_192_ _093_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ clknet_2_3__leaf_scan_clk _021_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_244_ clknet_2_0__leaf_scan_clk _006_ net5 VGND VGND VPWR VPWR GTC.col_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_175_ TIER1.MSS.scan_chain\[7\] _061_ _081_ TIER1.PRAS.scan_out VGND VGND VPWR VPWR
+ _082_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ net2 net26 _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ net58 net56 _108_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__mux2_1
Xhold6 GTC.shift_en VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ clknet_2_3__leaf_scan_clk _020_ net9 VGND VGND VPWR VPWR TIER1.MSS.scan_chain\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_191_ net37 net53 _091_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_243_ clknet_2_0__leaf_scan_clk _005_ net5 VGND VGND VPWR VPWR GTC.cluster_sel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_174_ GTC.mode_sel\[1\] GTC.mode_sel\[0\] VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__or2b_1
X_157_ _052_ _062_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_4
X_226_ net30 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__clkbuf_1
Xhold7 GTC.col_addr\[3\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_209_ _065_ GTC.mode_sel\[0\] _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_190_ _092_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_173_ net41 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
X_242_ clknet_2_0__leaf_scan_clk _004_ net5 VGND VGND VPWR VPWR GTC.cluster_sel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_156_ _071_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__clkbuf_1
X_225_ net29 TIER3.MSS.scan_chain\[4\] _108_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__mux2_1
Xhold8 GTC.tier_sel\[1\] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
X_208_ net3 GTC.tier_sel\[2\] VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2_1
X_139_ net25 _057_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_172_ net40 TIER1.MSS.scan_chain\[7\] _072_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__mux2_1
X_241_ clknet_2_0__leaf_scan_clk _003_ net5 VGND VGND VPWR VPWR GTC.shift_en sky130_fd_sc_hd__dfrtp_1
X_155_ net61 _070_ _049_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__mux2_1
X_224_ _112_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 _001_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
X_138_ GTC.col_addr\[2\] _057_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__and2_1
X_207_ net11 _101_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_171_ net33 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
X_240_ clknet_2_0__leaf_scan_clk _002_ net5 VGND VGND VPWR VPWR GTC.capture_en sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_223_ net46 net29 _108_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_154_ GTC.misr_t2 GTC.misr_t1 GTC.misr_t3 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_137_ _057_ _058_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__nor2_1
X_206_ _065_ TIER2.LC.scan_out _051_ _100_ GTC.capture_en VGND VGND VPWR VPWR _101_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_24_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_170_ net32 TIER1.MSS.scan_chain\[6\] _072_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_299_ GTC.cluster_sel\[1\] VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__buf_2
XFILLER_0_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_222_ _111_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__clkbuf_1
X_153_ _069_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_136_ _049_ net20 net22 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a21oi_1
X_205_ TIER2.MSS.scan_chain\[7\] _061_ _081_ TIER2.PRAS.scan_out VGND VGND VPWR VPWR
+ _100_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ GTC.cluster_sel\[0\] VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_152_ net57 net2 _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__mux2_1
X_221_ net48 net46 _108_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__mux2_1
X_204_ net50 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net3 GTC.col_addr\[0\] GTC.col_addr\[1\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_297_ TIER1.tier_sel\[1\] VGND VGND VPWR VPWR _297_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_220_ _110_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__clkbuf_1
X_151_ GTC.mode_sel\[0\] _052_ GTC.mode_sel\[1\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and3b_1
X_203_ net49 TIER2.MSS.scan_chain\[7\] _091_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__mux2_1
X_134_ _049_ net20 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput4 net4 VGND VGND VPWR VPWR fault_flag sky130_fd_sc_hd__clkbuf_4
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ GTC.capture_en VGND VGND VPWR VPWR _296_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_150_ _067_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ clknet_2_3__leaf_scan_clk _039_ net10 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_202_ net36 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_1
X_133_ net13 _055_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout5 net7 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 TIER3.LC.scan_out VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_295_ GTC.mode_sel\[1\] VGND VGND VPWR VPWR _295_/X sky130_fd_sc_hd__buf_2
XFILLER_0_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_278_ clknet_2_3__leaf_scan_clk _038_ net10 VGND VGND VPWR VPWR TIER3.MSS.scan_chain\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_201_ net35 TIER2.MSS.scan_chain\[6\] _091_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_132_ _056_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6 net7 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold40 _099_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net4 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

