module top_3d_jscan (fault_flag,
    reset_n,
    scan_clk,
    scan_in,
    test_enable);
 output fault_flag;
 input reset_n;
 input scan_clk;
 input scan_in;
 input test_enable;

 wire \GTC.capture_en ;
 wire \GTC.cluster_sel[0] ;
 wire \GTC.cluster_sel[1] ;
 wire \GTC.col_addr[0] ;
 wire \GTC.col_addr[1] ;
 wire \GTC.col_addr[2] ;
 wire \GTC.col_addr[3] ;
 wire \GTC.misr_t1 ;
 wire \GTC.misr_t2 ;
 wire \GTC.misr_t3 ;
 wire \GTC.mode_sel[0] ;
 wire \GTC.mode_sel[1] ;
 wire \GTC.shift_en ;
 wire \GTC.tier_sel[0] ;
 wire \GTC.tier_sel[1] ;
 wire \GTC.tier_sel[2] ;
 wire \TIER1.LC.scan_out ;
 wire \TIER1.MSS.scan_chain[0] ;
 wire \TIER1.MSS.scan_chain[1] ;
 wire \TIER1.MSS.scan_chain[2] ;
 wire \TIER1.MSS.scan_chain[3] ;
 wire \TIER1.MSS.scan_chain[4] ;
 wire \TIER1.MSS.scan_chain[5] ;
 wire \TIER1.MSS.scan_chain[6] ;
 wire \TIER1.MSS.scan_chain[7] ;
 wire \TIER1.PRAS.scan_out ;
 wire \TIER1.tier_sel[0] ;
 wire \TIER1.tier_sel[1] ;
 wire \TIER2.LC.scan_out ;
 wire \TIER2.MSS.scan_chain[0] ;
 wire \TIER2.MSS.scan_chain[1] ;
 wire \TIER2.MSS.scan_chain[2] ;
 wire \TIER2.MSS.scan_chain[3] ;
 wire \TIER2.MSS.scan_chain[4] ;
 wire \TIER2.MSS.scan_chain[5] ;
 wire \TIER2.MSS.scan_chain[6] ;
 wire \TIER2.MSS.scan_chain[7] ;
 wire \TIER2.PRAS.scan_out ;
 wire \TIER3.LC.scan_out ;
 wire \TIER3.MSS.scan_chain[0] ;
 wire \TIER3.MSS.scan_chain[1] ;
 wire \TIER3.MSS.scan_chain[2] ;
 wire \TIER3.MSS.scan_chain[3] ;
 wire \TIER3.MSS.scan_chain[4] ;
 wire \TIER3.MSS.scan_chain[5] ;
 wire \TIER3.MSS.scan_chain[6] ;
 wire \TIER3.MSS.scan_chain[7] ;
 wire \TIER3.PRAS.scan_out ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire capture_en;
 wire \cluster_sel[0] ;
 wire \cluster_sel[1] ;
 wire \col_addr[0] ;
 wire \col_addr[1] ;
 wire \col_addr[2] ;
 wire \col_addr[3] ;
 wire \mode_sel[0] ;
 wire \mode_sel[1] ;
 wire shift_en;
 wire test_en;
 wire \tier_sel[0] ;
 wire \tier_sel[1] ;
 wire tsv_scan_in;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;

 sky130_fd_sc_hd__clkbuf_4 _120_ (.A(net3),
    .X(_049_));
 sky130_fd_sc_hd__inv_2 _121_ (.A(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__and2_2 _122_ (.A(net3),
    .B(\GTC.tier_sel[1] ),
    .X(_051_));
 sky130_fd_sc_hd__a211o_1 _123_ (.A1(_050_),
    .A2(\GTC.tier_sel[0] ),
    .B1(_051_),
    .C1(\GTC.tier_sel[2] ),
    .X(_000_));
 sky130_fd_sc_hd__and2_2 _124_ (.A(net3),
    .B(\GTC.tier_sel[0] ),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _125_ (.A1(_050_),
    .A2(\GTC.tier_sel[2] ),
    .B1(\GTC.tier_sel[1] ),
    .C1(_052_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _126_ (.A0(\GTC.capture_en ),
    .A1(\GTC.shift_en ),
    .S(_049_),
    .X(_053_));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(_053_),
    .X(_002_));
 sky130_fd_sc_hd__xor2_1 _128_ (.A(_049_),
    .B(\GTC.shift_en ),
    .X(_003_));
 sky130_fd_sc_hd__or2_1 _129_ (.A(_049_),
    .B(\GTC.cluster_sel[0] ),
    .X(_054_));
 sky130_fd_sc_hd__nand2_1 _130_ (.A(_049_),
    .B(\GTC.cluster_sel[0] ),
    .Y(_055_));
 sky130_fd_sc_hd__and2_1 _131_ (.A(_054_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(_056_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _133_ (.A(\GTC.cluster_sel[1] ),
    .B(_055_),
    .Y(_005_));
 sky130_fd_sc_hd__xor2_1 _134_ (.A(_049_),
    .B(\GTC.col_addr[0] ),
    .X(_006_));
 sky130_fd_sc_hd__and3_1 _135_ (.A(net3),
    .B(\GTC.col_addr[0] ),
    .C(\GTC.col_addr[1] ),
    .X(_057_));
 sky130_fd_sc_hd__a21oi_1 _136_ (.A1(_049_),
    .A2(\GTC.col_addr[0] ),
    .B1(\GTC.col_addr[1] ),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _137_ (.A(_057_),
    .B(_058_),
    .Y(_007_));
 sky130_fd_sc_hd__and2_1 _138_ (.A(\GTC.col_addr[2] ),
    .B(_057_),
    .X(_059_));
 sky130_fd_sc_hd__nor2_1 _139_ (.A(\GTC.col_addr[2] ),
    .B(_057_),
    .Y(_060_));
 sky130_fd_sc_hd__nor2_1 _140_ (.A(_059_),
    .B(_060_),
    .Y(_008_));
 sky130_fd_sc_hd__xor2_1 _141_ (.A(\GTC.col_addr[3] ),
    .B(_059_),
    .X(_009_));
 sky130_fd_sc_hd__or2_2 _142_ (.A(\GTC.mode_sel[1] ),
    .B(\GTC.mode_sel[0] ),
    .X(_061_));
 sky130_fd_sc_hd__inv_2 _143_ (.A(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_1 _144_ (.A(\GTC.col_addr[3] ),
    .B(_059_),
    .Y(_063_));
 sky130_fd_sc_hd__mux2_1 _145_ (.A0(_062_),
    .A1(\GTC.mode_sel[0] ),
    .S(_063_),
    .X(_064_));
 sky130_fd_sc_hd__clkbuf_1 _146_ (.A(_064_),
    .X(_010_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(\GTC.mode_sel[1] ),
    .Y(_065_));
 sky130_fd_sc_hd__and2_1 _148_ (.A(_065_),
    .B(\GTC.mode_sel[0] ),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _149_ (.A0(_066_),
    .A1(\GTC.mode_sel[1] ),
    .S(_063_),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_1 _150_ (.A(_067_),
    .X(_011_));
 sky130_fd_sc_hd__and3b_1 _151_ (.A_N(\GTC.mode_sel[0] ),
    .B(_052_),
    .C(\GTC.mode_sel[1] ),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _152_ (.A0(\TIER1.LC.scan_out ),
    .A1(net2),
    .S(_068_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(_069_),
    .X(_012_));
 sky130_fd_sc_hd__or3_1 _154_ (.A(\GTC.misr_t2 ),
    .B(\GTC.misr_t1 ),
    .C(\GTC.misr_t3 ),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _155_ (.A0(net4),
    .A1(_070_),
    .S(_049_),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _156_ (.A(_071_),
    .X(_013_));
 sky130_fd_sc_hd__nand2_4 _157_ (.A(_052_),
    .B(_062_),
    .Y(_072_));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(net2),
    .A1(\TIER1.MSS.scan_chain[0] ),
    .S(_072_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _159_ (.A(_073_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(\TIER1.MSS.scan_chain[0] ),
    .A1(\TIER1.MSS.scan_chain[1] ),
    .S(_072_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(_074_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(\TIER1.MSS.scan_chain[1] ),
    .A1(\TIER1.MSS.scan_chain[2] ),
    .S(_072_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _163_ (.A(_075_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(\TIER1.MSS.scan_chain[2] ),
    .A1(\TIER1.MSS.scan_chain[3] ),
    .S(_072_),
    .X(_076_));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(_076_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _166_ (.A0(\TIER1.MSS.scan_chain[3] ),
    .A1(\TIER1.MSS.scan_chain[4] ),
    .S(_072_),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_1 _167_ (.A(_077_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\TIER1.MSS.scan_chain[4] ),
    .A1(\TIER1.MSS.scan_chain[5] ),
    .S(_072_),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(_078_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _170_ (.A0(\TIER1.MSS.scan_chain[5] ),
    .A1(\TIER1.MSS.scan_chain[6] ),
    .S(_072_),
    .X(_079_));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(_079_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(\TIER1.MSS.scan_chain[6] ),
    .A1(\TIER1.MSS.scan_chain[7] ),
    .S(_072_),
    .X(_080_));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(_080_),
    .X(_021_));
 sky130_fd_sc_hd__or2b_1 _174_ (.A(\GTC.mode_sel[1] ),
    .B_N(\GTC.mode_sel[0] ),
    .X(_081_));
 sky130_fd_sc_hd__o22a_1 _175_ (.A1(\TIER1.MSS.scan_chain[7] ),
    .A2(_061_),
    .B1(_081_),
    .B2(\TIER1.PRAS.scan_out ),
    .X(_082_));
 sky130_fd_sc_hd__o2111a_1 _176_ (.A1(_065_),
    .A2(\TIER1.LC.scan_out ),
    .B1(_052_),
    .C1(_082_),
    .D1(\GTC.capture_en ),
    .X(_083_));
 sky130_fd_sc_hd__xor2_1 _177_ (.A(\GTC.misr_t1 ),
    .B(_083_),
    .X(_022_));
 sky130_fd_sc_hd__xnor2_1 _178_ (.A(\GTC.col_addr[0] ),
    .B(\GTC.col_addr[2] ),
    .Y(_084_));
 sky130_fd_sc_hd__and4_1 _179_ (.A(_049_),
    .B(\GTC.tier_sel[2] ),
    .C(net8),
    .D(_066_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(\TIER3.PRAS.scan_out ),
    .A1(_084_),
    .S(_085_),
    .X(_086_));
 sky130_fd_sc_hd__clkbuf_1 _181_ (.A(_086_),
    .X(_023_));
 sky130_fd_sc_hd__and3b_1 _182_ (.A_N(\GTC.mode_sel[0] ),
    .B(_051_),
    .C(\GTC.mode_sel[1] ),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _183_ (.A0(\TIER2.LC.scan_out ),
    .A1(net2),
    .S(_087_),
    .X(_088_));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(_088_),
    .X(_024_));
 sky130_fd_sc_hd__and3_1 _185_ (.A(net8),
    .B(_052_),
    .C(_066_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _186_ (.A0(\TIER1.PRAS.scan_out ),
    .A1(_084_),
    .S(_089_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _187_ (.A(_090_),
    .X(_025_));
 sky130_fd_sc_hd__nand2_4 _188_ (.A(_051_),
    .B(_062_),
    .Y(_091_));
 sky130_fd_sc_hd__mux2_1 _189_ (.A0(net2),
    .A1(\TIER2.MSS.scan_chain[0] ),
    .S(_091_),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(_092_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _191_ (.A0(\TIER2.MSS.scan_chain[0] ),
    .A1(\TIER2.MSS.scan_chain[1] ),
    .S(_091_),
    .X(_093_));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(_093_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _193_ (.A0(\TIER2.MSS.scan_chain[1] ),
    .A1(\TIER2.MSS.scan_chain[2] ),
    .S(_091_),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(_094_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _195_ (.A0(\TIER2.MSS.scan_chain[2] ),
    .A1(\TIER2.MSS.scan_chain[3] ),
    .S(_091_),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(_095_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _197_ (.A0(\TIER2.MSS.scan_chain[3] ),
    .A1(\TIER2.MSS.scan_chain[4] ),
    .S(_091_),
    .X(_096_));
 sky130_fd_sc_hd__clkbuf_1 _198_ (.A(_096_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _199_ (.A0(\TIER2.MSS.scan_chain[4] ),
    .A1(\TIER2.MSS.scan_chain[5] ),
    .S(_091_),
    .X(_097_));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(_097_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _201_ (.A0(\TIER2.MSS.scan_chain[5] ),
    .A1(\TIER2.MSS.scan_chain[6] ),
    .S(_091_),
    .X(_098_));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(_098_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _203_ (.A0(\TIER2.MSS.scan_chain[6] ),
    .A1(\TIER2.MSS.scan_chain[7] ),
    .S(_091_),
    .X(_099_));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(_099_),
    .X(_033_));
 sky130_fd_sc_hd__o22a_1 _205_ (.A1(\TIER2.MSS.scan_chain[7] ),
    .A2(_061_),
    .B1(_081_),
    .B2(\TIER2.PRAS.scan_out ),
    .X(_100_));
 sky130_fd_sc_hd__o2111a_1 _206_ (.A1(_065_),
    .A2(\TIER2.LC.scan_out ),
    .B1(_051_),
    .C1(_100_),
    .D1(\GTC.capture_en ),
    .X(_101_));
 sky130_fd_sc_hd__xor2_1 _207_ (.A(\GTC.misr_t2 ),
    .B(_101_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _208_ (.A(net3),
    .B(\GTC.tier_sel[2] ),
    .Y(_102_));
 sky130_fd_sc_hd__or3_1 _209_ (.A(_065_),
    .B(\GTC.mode_sel[0] ),
    .C(_102_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _210_ (.A0(net2),
    .A1(\TIER3.LC.scan_out ),
    .S(_103_),
    .X(_104_));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(_104_),
    .X(_035_));
 sky130_fd_sc_hd__and3_1 _212_ (.A(net5),
    .B(_051_),
    .C(_066_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _213_ (.A0(\TIER2.PRAS.scan_out ),
    .A1(_084_),
    .S(_105_),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_1 _214_ (.A(_106_),
    .X(_036_));
 sky130_fd_sc_hd__or2_1 _215_ (.A(_061_),
    .B(_102_),
    .X(_107_));
 sky130_fd_sc_hd__buf_2 _216_ (.A(_107_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _217_ (.A0(net2),
    .A1(\TIER3.MSS.scan_chain[0] ),
    .S(_108_),
    .X(_109_));
 sky130_fd_sc_hd__clkbuf_1 _218_ (.A(_109_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _219_ (.A0(\TIER3.MSS.scan_chain[0] ),
    .A1(\TIER3.MSS.scan_chain[1] ),
    .S(_108_),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_1 _220_ (.A(_110_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(\TIER3.MSS.scan_chain[1] ),
    .A1(\TIER3.MSS.scan_chain[2] ),
    .S(_108_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _222_ (.A(_111_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _223_ (.A0(\TIER3.MSS.scan_chain[2] ),
    .A1(\TIER3.MSS.scan_chain[3] ),
    .S(_108_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _224_ (.A(_112_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _225_ (.A0(\TIER3.MSS.scan_chain[3] ),
    .A1(\TIER3.MSS.scan_chain[4] ),
    .S(_108_),
    .X(_113_));
 sky130_fd_sc_hd__clkbuf_1 _226_ (.A(_113_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _227_ (.A0(\TIER3.MSS.scan_chain[4] ),
    .A1(\TIER3.MSS.scan_chain[5] ),
    .S(_108_),
    .X(_114_));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(_114_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _229_ (.A0(\TIER3.MSS.scan_chain[5] ),
    .A1(\TIER3.MSS.scan_chain[6] ),
    .S(_108_),
    .X(_115_));
 sky130_fd_sc_hd__clkbuf_1 _230_ (.A(_115_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _231_ (.A0(\TIER3.MSS.scan_chain[6] ),
    .A1(\TIER3.MSS.scan_chain[7] ),
    .S(_108_),
    .X(_116_));
 sky130_fd_sc_hd__clkbuf_1 _232_ (.A(_116_),
    .X(_044_));
 sky130_fd_sc_hd__and3_1 _233_ (.A(_049_),
    .B(\GTC.tier_sel[2] ),
    .C(\GTC.capture_en ),
    .X(_117_));
 sky130_fd_sc_hd__o22a_1 _234_ (.A1(\TIER3.MSS.scan_chain[7] ),
    .A2(_061_),
    .B1(_081_),
    .B2(\TIER3.PRAS.scan_out ),
    .X(_118_));
 sky130_fd_sc_hd__o211a_1 _235_ (.A1(_065_),
    .A2(\TIER3.LC.scan_out ),
    .B1(_117_),
    .C1(_118_),
    .X(_119_));
 sky130_fd_sc_hd__xor2_1 _236_ (.A(\GTC.misr_t3 ),
    .B(_119_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_1 _237_ (.A1(_050_),
    .A2(\GTC.tier_sel[2] ),
    .B1(_051_),
    .X(_046_));
 sky130_fd_sc_hd__a21o_1 _238_ (.A1(_050_),
    .A2(\GTC.tier_sel[1] ),
    .B1(_052_),
    .X(_047_));
 sky130_fd_sc_hd__a21bo_1 _239_ (.A1(_050_),
    .A2(\GTC.tier_sel[0] ),
    .B1_N(_102_),
    .X(_048_));
 sky130_fd_sc_hd__dfrtp_1 _240_ (.CLK(scan_clk),
    .D(_002_),
    .RESET_B(net5),
    .Q(\GTC.capture_en ));
 sky130_fd_sc_hd__dfrtp_1 _241_ (.CLK(scan_clk),
    .D(_003_),
    .RESET_B(net5),
    .Q(\GTC.shift_en ));
 sky130_fd_sc_hd__dfrtp_1 _242_ (.CLK(scan_clk),
    .D(_004_),
    .RESET_B(net5),
    .Q(\GTC.cluster_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _243_ (.CLK(scan_clk),
    .D(_005_),
    .RESET_B(net5),
    .Q(\GTC.cluster_sel[1] ));
 sky130_fd_sc_hd__dfrtp_2 _244_ (.CLK(scan_clk),
    .D(_006_),
    .RESET_B(net5),
    .Q(\GTC.col_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _245_ (.CLK(scan_clk),
    .D(_007_),
    .RESET_B(net5),
    .Q(\GTC.col_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _246_ (.CLK(scan_clk),
    .D(_008_),
    .RESET_B(net5),
    .Q(\GTC.col_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _247_ (.CLK(scan_clk),
    .D(_009_),
    .RESET_B(net5),
    .Q(\GTC.col_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _248_ (.CLK(scan_clk),
    .D(_010_),
    .RESET_B(net6),
    .Q(\GTC.mode_sel[0] ));
 sky130_fd_sc_hd__dfrtp_2 _249_ (.CLK(scan_clk),
    .D(_011_),
    .RESET_B(net7),
    .Q(\GTC.mode_sel[1] ));
 sky130_fd_sc_hd__dfstp_1 _250_ (.CLK(scan_clk),
    .D(_000_),
    .SET_B(net8),
    .Q(\TIER1.tier_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _251_ (.CLK(scan_clk),
    .D(_001_),
    .RESET_B(net8),
    .Q(\TIER1.tier_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _252_ (.CLK(scan_clk),
    .D(_012_),
    .RESET_B(net9),
    .Q(\TIER1.LC.scan_out ));
 sky130_fd_sc_hd__dfrtp_1 _253_ (.CLK(scan_clk),
    .D(_013_),
    .RESET_B(net6),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _254_ (.CLK(scan_clk),
    .D(_014_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _255_ (.CLK(scan_clk),
    .D(_015_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[1] ));
 sky130_fd_sc_hd__dfrtp_1 _256_ (.CLK(scan_clk),
    .D(_016_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[2] ));
 sky130_fd_sc_hd__dfrtp_1 _257_ (.CLK(scan_clk),
    .D(_017_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[3] ));
 sky130_fd_sc_hd__dfrtp_1 _258_ (.CLK(scan_clk),
    .D(_018_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[4] ));
 sky130_fd_sc_hd__dfrtp_1 _259_ (.CLK(scan_clk),
    .D(_019_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[5] ));
 sky130_fd_sc_hd__dfrtp_1 _260_ (.CLK(scan_clk),
    .D(_020_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[6] ));
 sky130_fd_sc_hd__dfrtp_1 _261_ (.CLK(scan_clk),
    .D(_021_),
    .RESET_B(net9),
    .Q(\TIER1.MSS.scan_chain[7] ));
 sky130_fd_sc_hd__dfrtp_1 _262_ (.CLK(scan_clk),
    .D(_022_),
    .RESET_B(net6),
    .Q(\GTC.misr_t1 ));
 sky130_fd_sc_hd__dfxtp_1 _263_ (.CLK(scan_clk),
    .D(_023_),
    .Q(\TIER3.PRAS.scan_out ));
 sky130_fd_sc_hd__dfrtp_1 _264_ (.CLK(scan_clk),
    .D(_024_),
    .RESET_B(net6),
    .Q(\TIER2.LC.scan_out ));
 sky130_fd_sc_hd__dfxtp_1 _265_ (.CLK(scan_clk),
    .D(_025_),
    .Q(\TIER1.PRAS.scan_out ));
 sky130_fd_sc_hd__dfrtp_1 _266_ (.CLK(scan_clk),
    .D(_026_),
    .RESET_B(net6),
    .Q(\TIER2.MSS.scan_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _267_ (.CLK(scan_clk),
    .D(_027_),
    .RESET_B(net7),
    .Q(\TIER2.MSS.scan_chain[1] ));
 sky130_fd_sc_hd__dfrtp_1 _268_ (.CLK(scan_clk),
    .D(_028_),
    .RESET_B(net7),
    .Q(\TIER2.MSS.scan_chain[2] ));
 sky130_fd_sc_hd__dfrtp_1 _269_ (.CLK(scan_clk),
    .D(_029_),
    .RESET_B(net6),
    .Q(\TIER2.MSS.scan_chain[3] ));
 sky130_fd_sc_hd__dfrtp_1 _270_ (.CLK(scan_clk),
    .D(_030_),
    .RESET_B(net6),
    .Q(\TIER2.MSS.scan_chain[4] ));
 sky130_fd_sc_hd__dfrtp_1 _271_ (.CLK(scan_clk),
    .D(_031_),
    .RESET_B(net6),
    .Q(\TIER2.MSS.scan_chain[5] ));
 sky130_fd_sc_hd__dfrtp_1 _272_ (.CLK(scan_clk),
    .D(_032_),
    .RESET_B(net6),
    .Q(\TIER2.MSS.scan_chain[6] ));
 sky130_fd_sc_hd__dfrtp_1 _273_ (.CLK(scan_clk),
    .D(_033_),
    .RESET_B(net7),
    .Q(\TIER2.MSS.scan_chain[7] ));
 sky130_fd_sc_hd__dfrtp_1 _274_ (.CLK(scan_clk),
    .D(_034_),
    .RESET_B(net6),
    .Q(\GTC.misr_t2 ));
 sky130_fd_sc_hd__dfrtp_1 _275_ (.CLK(scan_clk),
    .D(_035_),
    .RESET_B(net9),
    .Q(\TIER3.LC.scan_out ));
 sky130_fd_sc_hd__dfxtp_1 _276_ (.CLK(scan_clk),
    .D(_036_),
    .Q(\TIER2.PRAS.scan_out ));
 sky130_fd_sc_hd__dfrtp_1 _277_ (.CLK(scan_clk),
    .D(_037_),
    .RESET_B(net10),
    .Q(\TIER3.MSS.scan_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _278_ (.CLK(scan_clk),
    .D(_038_),
    .RESET_B(net10),
    .Q(\TIER3.MSS.scan_chain[1] ));
 sky130_fd_sc_hd__dfrtp_1 _279_ (.CLK(scan_clk),
    .D(_039_),
    .RESET_B(net10),
    .Q(\TIER3.MSS.scan_chain[2] ));
 sky130_fd_sc_hd__dfrtp_1 _280_ (.CLK(scan_clk),
    .D(_040_),
    .RESET_B(net10),
    .Q(\TIER3.MSS.scan_chain[3] ));
 sky130_fd_sc_hd__dfrtp_1 _281_ (.CLK(scan_clk),
    .D(_041_),
    .RESET_B(net8),
    .Q(\TIER3.MSS.scan_chain[4] ));
 sky130_fd_sc_hd__dfrtp_1 _282_ (.CLK(scan_clk),
    .D(_042_),
    .RESET_B(net8),
    .Q(\TIER3.MSS.scan_chain[5] ));
 sky130_fd_sc_hd__dfrtp_1 _283_ (.CLK(scan_clk),
    .D(_043_),
    .RESET_B(net8),
    .Q(\TIER3.MSS.scan_chain[6] ));
 sky130_fd_sc_hd__dfrtp_1 _284_ (.CLK(scan_clk),
    .D(_044_),
    .RESET_B(net10),
    .Q(\TIER3.MSS.scan_chain[7] ));
 sky130_fd_sc_hd__dfrtp_1 _285_ (.CLK(scan_clk),
    .D(_045_),
    .RESET_B(net5),
    .Q(\GTC.misr_t3 ));
 sky130_fd_sc_hd__dfrtp_1 _286_ (.CLK(scan_clk),
    .D(_046_),
    .RESET_B(net8),
    .Q(\GTC.tier_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _287_ (.CLK(scan_clk),
    .D(_047_),
    .RESET_B(net8),
    .Q(\GTC.tier_sel[1] ));
 sky130_fd_sc_hd__dfstp_1 _288_ (.CLK(scan_clk),
    .D(_048_),
    .SET_B(net8),
    .Q(\GTC.tier_sel[0] ));
 sky130_fd_sc_hd__buf_2 _289_ (.A(\GTC.col_addr[0] ),
    .X(\col_addr[0] ));
 sky130_fd_sc_hd__buf_2 _290_ (.A(\TIER1.tier_sel[0] ),
    .X(\tier_sel[0] ));
 sky130_fd_sc_hd__buf_2 _291_ (.A(\GTC.col_addr[1] ),
    .X(\col_addr[1] ));
 sky130_fd_sc_hd__buf_2 _292_ (.A(\GTC.col_addr[2] ),
    .X(\col_addr[2] ));
 sky130_fd_sc_hd__buf_2 _293_ (.A(\GTC.col_addr[3] ),
    .X(\col_addr[3] ));
 sky130_fd_sc_hd__buf_2 _294_ (.A(\GTC.mode_sel[0] ),
    .X(\mode_sel[0] ));
 sky130_fd_sc_hd__buf_2 _295_ (.A(\GTC.mode_sel[1] ),
    .X(\mode_sel[1] ));
 sky130_fd_sc_hd__buf_2 _296_ (.A(\GTC.capture_en ),
    .X(capture_en));
 sky130_fd_sc_hd__buf_2 _297_ (.A(\TIER1.tier_sel[1] ),
    .X(\tier_sel[1] ));
 sky130_fd_sc_hd__buf_2 _298_ (.A(\GTC.cluster_sel[0] ),
    .X(\cluster_sel[0] ));
 sky130_fd_sc_hd__buf_2 _299_ (.A(\GTC.cluster_sel[1] ),
    .X(\cluster_sel[1] ));
 sky130_fd_sc_hd__buf_2 _300_ (.A(\GTC.shift_en ),
    .X(shift_en));
 sky130_fd_sc_hd__buf_2 _301_ (.A(net3),
    .X(test_en));
 sky130_fd_sc_hd__buf_2 _302_ (.A(net2),
    .X(tsv_scan_in));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(reset_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(scan_in),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(test_enable),
    .X(net3));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(fault_flag));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net7),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 fanout6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 fanout7 (.A(net1),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net10),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net1),
    .X(net10));
endmodule
