magic
tech sky130A
magscale 1 2
timestamp 1772104682
<< obsli1 >>
rect 1104 2159 16284 16881
<< obsm1 >>
rect 14 2128 16284 16912
<< metal2 >>
rect 9678 18774 9734 19574
rect 18 0 74 800
rect 14186 0 14242 800
<< obsm2 >>
rect 20 18718 9622 18774
rect 9790 18718 15896 18774
rect 20 856 15896 18718
rect 130 800 14130 856
rect 14298 800 15896 856
<< metal3 >>
rect 0 14968 800 15088
rect 16630 11568 17430 11688
<< obsm3 >>
rect 798 15168 16630 16897
rect 880 14888 16630 15168
rect 798 11768 16630 14888
rect 798 11488 16550 11768
rect 798 2143 16630 11488
<< metal4 >>
rect 2841 2128 3161 16912
rect 3501 2128 3821 16912
rect 6636 2128 6956 16912
rect 7296 2128 7616 16912
rect 10431 2128 10751 16912
rect 11091 2128 11411 16912
rect 14226 2128 14546 16912
rect 14886 2128 15206 16912
<< obsm4 >>
rect 13675 9555 13741 11661
<< metal5 >>
rect 1056 15528 16332 15848
rect 1056 14868 16332 15188
rect 1056 11856 16332 12176
rect 1056 11196 16332 11516
rect 1056 8184 16332 8504
rect 1056 7524 16332 7844
rect 1056 4512 16332 4832
rect 1056 3852 16332 4172
<< labels >>
rlabel metal4 s 3501 2128 3821 16912 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7296 2128 7616 16912 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11091 2128 11411 16912 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14886 2128 15206 16912 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4512 16332 4832 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8184 16332 8504 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11856 16332 12176 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 15528 16332 15848 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2841 2128 3161 16912 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6636 2128 6956 16912 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10431 2128 10751 16912 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14226 2128 14546 16912 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3852 16332 4172 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7524 16332 7844 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11196 16332 11516 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 14868 16332 15188 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 14968 800 15088 6 fault_flag
port 3 nsew signal output
rlabel metal2 s 18 0 74 800 6 reset_n
port 4 nsew signal input
rlabel metal3 s 16630 11568 17430 11688 6 scan_clk
port 5 nsew signal input
rlabel metal2 s 9678 18774 9734 19574 6 scan_in
port 6 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 test_enable
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 17430 19574
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 837758
string GDS_FILE /openlane/designs/jscan/runs/RUN_2026.02.26_11.15.28/results/signoff/top_3d_jscan.magic.gds
string GDS_START 260046
<< end >>

