magic
tech sky130A
magscale 1 2
timestamp 1772104692
<< checkpaint >>
rect -3932 -3932 21362 23506
<< viali >>
rect 10057 16609 10091 16643
rect 9873 16541 9907 16575
rect 6561 16065 6595 16099
rect 4537 15997 4571 16031
rect 5273 15997 5307 16031
rect 6745 15997 6779 16031
rect 7389 15997 7423 16031
rect 9597 15997 9631 16031
rect 9781 15997 9815 16031
rect 12081 15997 12115 16031
rect 3985 15861 4019 15895
rect 4721 15861 4755 15895
rect 6377 15861 6411 15895
rect 9045 15861 9079 15895
rect 10425 15861 10459 15895
rect 11529 15861 11563 15895
rect 6088 15657 6122 15691
rect 7573 15657 7607 15691
rect 9505 15657 9539 15691
rect 3893 15521 3927 15555
rect 5825 15521 5859 15555
rect 10057 15521 10091 15555
rect 10425 15521 10459 15555
rect 10609 15521 10643 15555
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 5549 15453 5583 15487
rect 8309 15453 8343 15487
rect 8677 15453 8711 15487
rect 9137 15453 9171 15487
rect 9413 15453 9447 15487
rect 9873 15453 9907 15487
rect 11161 15453 11195 15487
rect 11805 15453 11839 15487
rect 14657 15453 14691 15487
rect 1777 15385 1811 15419
rect 4077 15385 4111 15419
rect 5273 15385 5307 15419
rect 12081 15385 12115 15419
rect 1501 15317 1535 15351
rect 4537 15317 4571 15351
rect 5733 15317 5767 15351
rect 7665 15317 7699 15351
rect 8953 15317 8987 15351
rect 9229 15317 9263 15351
rect 9965 15317 9999 15351
rect 10701 15317 10735 15351
rect 11069 15317 11103 15351
rect 11345 15317 11379 15351
rect 13553 15317 13587 15351
rect 14105 15317 14139 15351
rect 4353 15113 4387 15147
rect 4445 15113 4479 15147
rect 7297 15113 7331 15147
rect 9505 15113 9539 15147
rect 11345 15113 11379 15147
rect 13277 15113 13311 15147
rect 13737 15113 13771 15147
rect 5917 15045 5951 15079
rect 8033 15045 8067 15079
rect 6193 14977 6227 15011
rect 6745 14977 6779 15011
rect 7205 14977 7239 15011
rect 7757 14977 7791 15011
rect 14749 14977 14783 15011
rect 2605 14909 2639 14943
rect 2881 14909 2915 14943
rect 7389 14909 7423 14943
rect 9597 14909 9631 14943
rect 9873 14909 9907 14943
rect 11529 14909 11563 14943
rect 11805 14909 11839 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 6837 14841 6871 14875
rect 14197 14841 14231 14875
rect 6561 14773 6595 14807
rect 13369 14773 13403 14807
rect 3893 14569 3927 14603
rect 5365 14569 5399 14603
rect 7941 14569 7975 14603
rect 10793 14569 10827 14603
rect 3617 14501 3651 14535
rect 10701 14501 10735 14535
rect 1869 14433 1903 14467
rect 4537 14433 4571 14467
rect 5917 14433 5951 14467
rect 6469 14433 6503 14467
rect 8953 14433 8987 14467
rect 11253 14433 11287 14467
rect 13921 14433 13955 14467
rect 4077 14365 4111 14399
rect 4353 14365 4387 14399
rect 4813 14365 4847 14399
rect 6193 14365 6227 14399
rect 10977 14365 11011 14399
rect 2145 14297 2179 14331
rect 9229 14297 9263 14331
rect 13645 14297 13679 14331
rect 4169 14229 4203 14263
rect 4721 14229 4755 14263
rect 5181 14229 5215 14263
rect 5733 14229 5767 14263
rect 5825 14229 5859 14263
rect 11437 14229 11471 14263
rect 11529 14229 11563 14263
rect 11897 14229 11931 14263
rect 12173 14229 12207 14263
rect 4261 14025 4295 14059
rect 4721 14025 4755 14059
rect 6561 14025 6595 14059
rect 6929 14025 6963 14059
rect 9229 14025 9263 14059
rect 9689 14025 9723 14059
rect 10701 14025 10735 14059
rect 11529 14025 11563 14059
rect 13185 14025 13219 14059
rect 14013 14025 14047 14059
rect 2789 13957 2823 13991
rect 7021 13957 7055 13991
rect 12725 13957 12759 13991
rect 12817 13957 12851 13991
rect 4813 13889 4847 13923
rect 5181 13889 5215 13923
rect 5733 13889 5767 13923
rect 9597 13889 9631 13923
rect 11253 13889 11287 13923
rect 12081 13889 12115 13923
rect 14197 13889 14231 13923
rect 2513 13821 2547 13855
rect 4997 13821 5031 13855
rect 7113 13821 7147 13855
rect 9781 13821 9815 13855
rect 12633 13821 12667 13855
rect 13829 13821 13863 13855
rect 13277 13753 13311 13787
rect 4353 13685 4387 13719
rect 3065 13481 3099 13515
rect 11805 13481 11839 13515
rect 12909 13413 12943 13447
rect 5089 13345 5123 13379
rect 5825 13345 5859 13379
rect 12357 13345 12391 13379
rect 13553 13345 13587 13379
rect 3249 13277 3283 13311
rect 4813 13277 4847 13311
rect 6561 13277 6595 13311
rect 7297 13277 7331 13311
rect 11621 13277 11655 13311
rect 12081 13277 12115 13311
rect 13001 13277 13035 13311
rect 4905 13209 4939 13243
rect 12541 13209 12575 13243
rect 4445 13141 4479 13175
rect 5273 13141 5307 13175
rect 6009 13141 6043 13175
rect 6745 13141 6779 13175
rect 11897 13141 11931 13175
rect 12449 13141 12483 13175
rect 5825 12937 5859 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 13277 12937 13311 12971
rect 11805 12869 11839 12903
rect 6837 12801 6871 12835
rect 11529 12801 11563 12835
rect 13921 12801 13955 12835
rect 4077 12733 4111 12767
rect 4353 12733 4387 12767
rect 7021 12733 7055 12767
rect 13369 12597 13403 12631
rect 4261 12393 4295 12427
rect 11437 12325 11471 12359
rect 2237 12257 2271 12291
rect 5089 12257 5123 12291
rect 5825 12257 5859 12291
rect 7573 12257 7607 12291
rect 11345 12257 11379 12291
rect 11989 12257 12023 12291
rect 3157 12189 3191 12223
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 5549 12189 5583 12223
rect 8217 12189 8251 12223
rect 9781 12189 9815 12223
rect 11805 12189 11839 12223
rect 14657 12189 14691 12223
rect 15025 12189 15059 12223
rect 15853 12189 15887 12223
rect 6101 12121 6135 12155
rect 2881 12053 2915 12087
rect 2973 12053 3007 12087
rect 5733 12053 5767 12087
rect 7665 12053 7699 12087
rect 9229 12053 9263 12087
rect 10701 12053 10735 12087
rect 11897 12053 11931 12087
rect 14105 12053 14139 12087
rect 14841 12053 14875 12087
rect 15301 12053 15335 12087
rect 1501 11849 1535 11883
rect 6929 11849 6963 11883
rect 7297 11849 7331 11883
rect 7389 11849 7423 11883
rect 12817 11849 12851 11883
rect 14657 11849 14691 11883
rect 14749 11849 14783 11883
rect 10517 11781 10551 11815
rect 13185 11781 13219 11815
rect 6653 11713 6687 11747
rect 11253 11713 11287 11747
rect 12633 11713 12667 11747
rect 15117 11713 15151 11747
rect 2973 11645 3007 11679
rect 3249 11645 3283 11679
rect 7481 11645 7515 11679
rect 8309 11645 8343 11679
rect 8585 11645 8619 11679
rect 12909 11645 12943 11679
rect 15209 11645 15243 11679
rect 15393 11645 15427 11679
rect 6469 11509 6503 11543
rect 10057 11509 10091 11543
rect 10241 11509 10275 11543
rect 11069 11509 11103 11543
rect 3249 11305 3283 11339
rect 6088 11305 6122 11339
rect 7573 11305 7607 11339
rect 8953 11305 8987 11339
rect 10780 11305 10814 11339
rect 13093 11305 13127 11339
rect 14368 11305 14402 11339
rect 15853 11305 15887 11339
rect 8769 11237 8803 11271
rect 13001 11237 13035 11271
rect 2697 11169 2731 11203
rect 5825 11169 5859 11203
rect 8217 11169 8251 11203
rect 9689 11169 9723 11203
rect 10517 11169 10551 11203
rect 12265 11169 12299 11203
rect 13553 11169 13587 11203
rect 13645 11169 13679 11203
rect 2881 11101 2915 11135
rect 8401 11101 8435 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9873 11101 9907 11135
rect 10149 11101 10183 11135
rect 12817 11101 12851 11135
rect 13461 11101 13495 11135
rect 14105 11101 14139 11135
rect 2789 10965 2823 10999
rect 8309 10965 8343 10999
rect 10333 10965 10367 10999
rect 7205 10761 7239 10795
rect 4537 10693 4571 10727
rect 7021 10693 7055 10727
rect 11069 10693 11103 10727
rect 13829 10693 13863 10727
rect 2237 10625 2271 10659
rect 4169 10625 4203 10659
rect 7297 10625 7331 10659
rect 7665 10625 7699 10659
rect 8033 10625 8067 10659
rect 8401 10625 8435 10659
rect 8769 10625 8803 10659
rect 11345 10625 11379 10659
rect 13553 10625 13587 10659
rect 2513 10557 2547 10591
rect 8953 10557 8987 10591
rect 6653 10489 6687 10523
rect 3985 10421 4019 10455
rect 7021 10421 7055 10455
rect 9505 10421 9539 10455
rect 9597 10421 9631 10455
rect 15301 10421 15335 10455
rect 2145 10217 2179 10251
rect 2237 10217 2271 10251
rect 5733 10217 5767 10251
rect 7757 10217 7791 10251
rect 8953 10217 8987 10251
rect 9137 10217 9171 10251
rect 10333 10217 10367 10251
rect 11897 10217 11931 10251
rect 14289 10217 14323 10251
rect 8033 10149 8067 10183
rect 15117 10149 15151 10183
rect 2697 10081 2731 10115
rect 3525 10081 3559 10115
rect 4537 10081 4571 10115
rect 4997 10081 5031 10115
rect 7113 10081 7147 10115
rect 8677 10081 8711 10115
rect 9781 10081 9815 10115
rect 9873 10081 9907 10115
rect 14933 10081 14967 10115
rect 15669 10081 15703 10115
rect 2053 10013 2087 10047
rect 2145 10013 2179 10047
rect 2605 10013 2639 10047
rect 2881 10013 2915 10047
rect 3893 10013 3927 10047
rect 4445 10013 4479 10047
rect 4905 10013 4939 10047
rect 7389 10013 7423 10047
rect 7481 10013 7515 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 8769 10013 8803 10047
rect 9505 10013 9539 10047
rect 10425 10013 10459 10047
rect 14657 10013 14691 10047
rect 7021 9945 7055 9979
rect 8401 9945 8435 9979
rect 1777 9877 1811 9911
rect 7573 9877 7607 9911
rect 8493 9877 8527 9911
rect 9137 9877 9171 9911
rect 9965 9877 9999 9911
rect 14749 9877 14783 9911
rect 15485 9877 15519 9911
rect 15577 9877 15611 9911
rect 2421 9673 2455 9707
rect 7481 9673 7515 9707
rect 10609 9673 10643 9707
rect 15945 9673 15979 9707
rect 3893 9605 3927 9639
rect 6745 9605 6779 9639
rect 8953 9605 8987 9639
rect 5365 9537 5399 9571
rect 6101 9537 6135 9571
rect 6837 9537 6871 9571
rect 7665 9537 7699 9571
rect 7757 9537 7791 9571
rect 8033 9537 8067 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 10517 9537 10551 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11161 9537 11195 9571
rect 13185 9537 13219 9571
rect 15301 9537 15335 9571
rect 4169 9469 4203 9503
rect 4905 9469 4939 9503
rect 4997 9469 5031 9503
rect 5457 9469 5491 9503
rect 7021 9469 7055 9503
rect 7941 9469 7975 9503
rect 8309 9469 8343 9503
rect 13461 9469 13495 9503
rect 13737 9469 13771 9503
rect 6377 9401 6411 9435
rect 13369 9401 13403 9435
rect 4261 9333 4295 9367
rect 5917 9333 5951 9367
rect 11069 9333 11103 9367
rect 15209 9333 15243 9367
rect 1869 9129 1903 9163
rect 4445 9129 4479 9163
rect 8309 9129 8343 9163
rect 8677 9129 8711 9163
rect 9505 9129 9539 9163
rect 10609 9129 10643 9163
rect 10793 9129 10827 9163
rect 7389 9061 7423 9095
rect 12541 9061 12575 9095
rect 14841 9061 14875 9095
rect 3341 8993 3375 9027
rect 3801 8993 3835 9027
rect 5733 8993 5767 9027
rect 7941 8993 7975 9027
rect 9321 8993 9355 9027
rect 10885 8993 10919 9027
rect 14289 8993 14323 9027
rect 3617 8925 3651 8959
rect 5457 8925 5491 8959
rect 7849 8925 7883 8959
rect 8217 8925 8251 8959
rect 9137 8925 9171 8959
rect 9413 8925 9447 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10977 8925 11011 8959
rect 11069 8925 11103 8959
rect 11437 8925 11471 8959
rect 12357 8925 12391 8959
rect 13461 8925 13495 8959
rect 14473 8925 14507 8959
rect 15485 8925 15519 8959
rect 7757 8857 7791 8891
rect 9689 8857 9723 8891
rect 11253 8857 11287 8891
rect 14933 8857 14967 8891
rect 7205 8789 7239 8823
rect 8953 8789 8987 8823
rect 12909 8789 12943 8823
rect 14381 8789 14415 8823
rect 8125 8585 8159 8619
rect 9229 8585 9263 8619
rect 10149 8585 10183 8619
rect 10793 8585 10827 8619
rect 10961 8585 10995 8619
rect 13001 8585 13035 8619
rect 15669 8585 15703 8619
rect 11161 8517 11195 8551
rect 13369 8517 13403 8551
rect 6009 8449 6043 8483
rect 8953 8449 8987 8483
rect 9321 8449 9355 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10701 8449 10735 8483
rect 11713 8449 11747 8483
rect 11989 8449 12023 8483
rect 12909 8449 12943 8483
rect 13921 8449 13955 8483
rect 14565 8449 14599 8483
rect 15117 8449 15151 8483
rect 6377 8381 6411 8415
rect 6653 8381 6687 8415
rect 9965 8381 9999 8415
rect 10609 8381 10643 8415
rect 12357 8381 12391 8415
rect 13461 8381 13495 8415
rect 13645 8381 13679 8415
rect 14289 8381 14323 8415
rect 14473 8381 14507 8415
rect 6193 8313 6227 8347
rect 8401 8245 8435 8279
rect 9413 8245 9447 8279
rect 10977 8245 11011 8279
rect 11529 8245 11563 8279
rect 12173 8245 12207 8279
rect 14105 8245 14139 8279
rect 14933 8245 14967 8279
rect 8493 8041 8527 8075
rect 9229 8041 9263 8075
rect 10885 8041 10919 8075
rect 13737 8041 13771 8075
rect 15853 8041 15887 8075
rect 2697 7973 2731 8007
rect 3249 7905 3283 7939
rect 12265 7905 12299 7939
rect 14381 7905 14415 7939
rect 2605 7837 2639 7871
rect 3065 7837 3099 7871
rect 4077 7837 4111 7871
rect 7113 7837 7147 7871
rect 9505 7837 9539 7871
rect 11989 7837 12023 7871
rect 14105 7837 14139 7871
rect 5273 7769 5307 7803
rect 7021 7769 7055 7803
rect 7380 7769 7414 7803
rect 9045 7769 9079 7803
rect 9772 7769 9806 7803
rect 2421 7701 2455 7735
rect 3157 7701 3191 7735
rect 9245 7701 9279 7735
rect 9413 7701 9447 7735
rect 3893 7497 3927 7531
rect 6929 7497 6963 7531
rect 7599 7497 7633 7531
rect 7849 7497 7883 7531
rect 8217 7497 8251 7531
rect 9137 7497 9171 7531
rect 9597 7497 9631 7531
rect 12817 7497 12851 7531
rect 15025 7497 15059 7531
rect 2329 7429 2363 7463
rect 7389 7429 7423 7463
rect 10732 7429 10766 7463
rect 15117 7429 15151 7463
rect 1593 7361 1627 7395
rect 4629 7361 4663 7395
rect 6745 7361 6779 7395
rect 9045 7361 9079 7395
rect 10977 7361 11011 7395
rect 15669 7361 15703 7395
rect 1685 7293 1719 7327
rect 2053 7293 2087 7327
rect 3801 7293 3835 7327
rect 4445 7293 4479 7327
rect 8309 7293 8343 7327
rect 8401 7293 8435 7327
rect 8953 7293 8987 7327
rect 14289 7293 14323 7327
rect 14565 7293 14599 7327
rect 15209 7293 15243 7327
rect 7757 7225 7791 7259
rect 9505 7225 9539 7259
rect 1961 7157 1995 7191
rect 7573 7157 7607 7191
rect 14657 7157 14691 7191
rect 15485 7157 15519 7191
rect 2126 6953 2160 6987
rect 11253 6953 11287 6987
rect 13553 6953 13587 6987
rect 14368 6953 14402 6987
rect 6377 6817 6411 6851
rect 9781 6817 9815 6851
rect 11069 6817 11103 6851
rect 14105 6817 14139 6851
rect 1869 6749 1903 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 11437 6749 11471 6783
rect 13369 6749 13403 6783
rect 9965 6681 9999 6715
rect 10517 6681 10551 6715
rect 3617 6613 3651 6647
rect 9873 6613 9907 6647
rect 10333 6613 10367 6647
rect 15853 6613 15887 6647
rect 2697 6409 2731 6443
rect 9505 6409 9539 6443
rect 9873 6409 9907 6443
rect 15209 6409 15243 6443
rect 9689 6341 9723 6375
rect 10057 6341 10091 6375
rect 3341 6273 3375 6307
rect 7113 6273 7147 6307
rect 9781 6273 9815 6307
rect 10793 6273 10827 6307
rect 15761 6273 15795 6307
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 6193 6205 6227 6239
rect 6929 6205 6963 6239
rect 6377 6069 6411 6103
rect 10977 6069 11011 6103
rect 5181 5865 5215 5899
rect 11897 5865 11931 5899
rect 15301 5865 15335 5899
rect 7205 5797 7239 5831
rect 5641 5729 5675 5763
rect 6745 5729 6779 5763
rect 15853 5729 15887 5763
rect 5549 5661 5583 5695
rect 6837 5661 6871 5695
rect 9665 5671 9699 5705
rect 9771 5639 9805 5673
rect 9873 5661 9907 5695
rect 10057 5661 10091 5695
rect 10157 5661 10191 5695
rect 10425 5661 10459 5695
rect 9597 5525 9631 5559
rect 10333 5525 10367 5559
rect 5825 5321 5859 5355
rect 9597 5321 9631 5355
rect 2881 5253 2915 5287
rect 6469 5253 6503 5287
rect 11345 5253 11379 5287
rect 2697 5185 2731 5219
rect 5549 5185 5583 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 9413 5185 9447 5219
rect 9689 5185 9723 5219
rect 12081 5185 12115 5219
rect 12265 5185 12299 5219
rect 12357 5185 12391 5219
rect 12541 5185 12575 5219
rect 12633 5185 12667 5219
rect 6193 5117 6227 5151
rect 7389 5117 7423 5151
rect 9965 5117 9999 5151
rect 10057 5117 10091 5151
rect 10425 5117 10459 5151
rect 10793 5117 10827 5151
rect 3065 4981 3099 5015
rect 5733 4981 5767 5015
rect 9229 4981 9263 5015
rect 9781 4981 9815 5015
rect 11529 4981 11563 5015
rect 12817 4981 12851 5015
rect 3249 4777 3283 4811
rect 7021 4777 7055 4811
rect 7297 4777 7331 4811
rect 8677 4777 8711 4811
rect 10885 4777 10919 4811
rect 11240 4777 11274 4811
rect 2605 4641 2639 4675
rect 5273 4641 5307 4675
rect 5549 4641 5583 4675
rect 9137 4641 9171 4675
rect 10977 4641 11011 4675
rect 2237 4573 2271 4607
rect 2697 4573 2731 4607
rect 3801 4573 3835 4607
rect 4353 4573 4387 4607
rect 4537 4573 4571 4607
rect 7573 4573 7607 4607
rect 8585 4573 8619 4607
rect 8769 4573 8803 4607
rect 3341 4505 3375 4539
rect 7481 4505 7515 4539
rect 9413 4505 9447 4539
rect 2053 4437 2087 4471
rect 2329 4437 2363 4471
rect 4721 4437 4755 4471
rect 7113 4437 7147 4471
rect 7281 4437 7315 4471
rect 12725 4437 12759 4471
rect 3893 4233 3927 4267
rect 9045 4233 9079 4267
rect 2329 4165 2363 4199
rect 6193 4165 6227 4199
rect 7573 4165 7607 4199
rect 1777 4097 1811 4131
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 4077 4097 4111 4131
rect 4169 4097 4203 4131
rect 4353 4097 4387 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 5917 4097 5951 4131
rect 6009 4097 6043 4131
rect 7205 4097 7239 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 9229 4097 9263 4131
rect 9597 4097 9631 4131
rect 11529 4097 11563 4131
rect 13323 4097 13357 4131
rect 13461 4097 13495 4131
rect 1869 4029 1903 4063
rect 11897 4029 11931 4063
rect 3801 3961 3835 3995
rect 6193 3961 6227 3995
rect 5825 3893 5859 3927
rect 6561 3893 6595 3927
rect 8677 3893 8711 3927
rect 11023 3893 11057 3927
rect 3525 3689 3559 3723
rect 7573 3689 7607 3723
rect 11069 3689 11103 3723
rect 8401 3621 8435 3655
rect 11805 3621 11839 3655
rect 1777 3553 1811 3587
rect 5457 3553 5491 3587
rect 5733 3553 5767 3587
rect 6101 3553 6135 3587
rect 9229 3553 9263 3587
rect 9505 3553 9539 3587
rect 10977 3553 11011 3587
rect 11621 3553 11655 3587
rect 12449 3553 12483 3587
rect 4077 3485 4111 3519
rect 5365 3485 5399 3519
rect 5825 3485 5859 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 12633 3485 12667 3519
rect 13553 3485 13587 3519
rect 2053 3417 2087 3451
rect 8125 3145 8159 3179
rect 10701 3145 10735 3179
rect 11621 3145 11655 3179
rect 6653 3077 6687 3111
rect 10149 3077 10183 3111
rect 6377 3009 6411 3043
rect 10333 3009 10367 3043
rect 10977 3009 11011 3043
rect 11805 3009 11839 3043
rect 10517 2941 10551 2975
rect 11989 2941 12023 2975
rect 1593 2601 1627 2635
rect 14381 2465 14415 2499
rect 1409 2397 1443 2431
rect 14105 2397 14139 2431
<< metal1 >>
rect 1104 16890 16284 16912
rect 1104 16838 2847 16890
rect 2899 16838 2911 16890
rect 2963 16838 2975 16890
rect 3027 16838 3039 16890
rect 3091 16838 3103 16890
rect 3155 16838 6642 16890
rect 6694 16838 6706 16890
rect 6758 16838 6770 16890
rect 6822 16838 6834 16890
rect 6886 16838 6898 16890
rect 6950 16838 10437 16890
rect 10489 16838 10501 16890
rect 10553 16838 10565 16890
rect 10617 16838 10629 16890
rect 10681 16838 10693 16890
rect 10745 16838 14232 16890
rect 14284 16838 14296 16890
rect 14348 16838 14360 16890
rect 14412 16838 14424 16890
rect 14476 16838 14488 16890
rect 14540 16838 16284 16890
rect 1104 16816 16284 16838
rect 10045 16643 10103 16649
rect 10045 16609 10057 16643
rect 10091 16640 10103 16643
rect 10226 16640 10232 16652
rect 10091 16612 10232 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 1104 16346 16284 16368
rect 1104 16294 3507 16346
rect 3559 16294 3571 16346
rect 3623 16294 3635 16346
rect 3687 16294 3699 16346
rect 3751 16294 3763 16346
rect 3815 16294 7302 16346
rect 7354 16294 7366 16346
rect 7418 16294 7430 16346
rect 7482 16294 7494 16346
rect 7546 16294 7558 16346
rect 7610 16294 11097 16346
rect 11149 16294 11161 16346
rect 11213 16294 11225 16346
rect 11277 16294 11289 16346
rect 11341 16294 11353 16346
rect 11405 16294 14892 16346
rect 14944 16294 14956 16346
rect 15008 16294 15020 16346
rect 15072 16294 15084 16346
rect 15136 16294 15148 16346
rect 15200 16294 16284 16346
rect 1104 16272 16284 16294
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 6512 16068 6561 16096
rect 6512 16056 6518 16068
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4396 16000 4537 16028
rect 4396 15988 4402 16000
rect 4525 15997 4537 16000
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 5258 15988 5264 16040
rect 5316 15988 5322 16040
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 6420 16000 6745 16028
rect 6420 15988 6426 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 7374 15988 7380 16040
rect 7432 15988 7438 16040
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 9766 15988 9772 16040
rect 9824 15988 9830 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11664 16000 12081 16028
rect 11664 15988 11670 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 3970 15852 3976 15904
rect 4028 15852 4034 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 4798 15892 4804 15904
rect 4755 15864 4804 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 6236 15864 6377 15892
rect 6236 15852 6242 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 6365 15855 6423 15861
rect 9030 15852 9036 15904
rect 9088 15852 9094 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 9916 15864 10425 15892
rect 9916 15852 9922 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 11514 15852 11520 15904
rect 11572 15852 11578 15904
rect 1104 15802 16284 15824
rect 1104 15750 2847 15802
rect 2899 15750 2911 15802
rect 2963 15750 2975 15802
rect 3027 15750 3039 15802
rect 3091 15750 3103 15802
rect 3155 15750 6642 15802
rect 6694 15750 6706 15802
rect 6758 15750 6770 15802
rect 6822 15750 6834 15802
rect 6886 15750 6898 15802
rect 6950 15750 10437 15802
rect 10489 15750 10501 15802
rect 10553 15750 10565 15802
rect 10617 15750 10629 15802
rect 10681 15750 10693 15802
rect 10745 15750 14232 15802
rect 14284 15750 14296 15802
rect 14348 15750 14360 15802
rect 14412 15750 14424 15802
rect 14476 15750 14488 15802
rect 14540 15750 16284 15802
rect 1104 15728 16284 15750
rect 6076 15691 6134 15697
rect 6076 15657 6088 15691
rect 6122 15688 6134 15691
rect 6178 15688 6184 15700
rect 6122 15660 6184 15688
rect 6122 15657 6134 15660
rect 6076 15651 6134 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 7374 15648 7380 15700
rect 7432 15688 7438 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7432 15660 7573 15688
rect 7432 15648 7438 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 9030 15648 9036 15700
rect 9088 15648 9094 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9582 15688 9588 15700
rect 9539 15660 9588 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15552 3939 15555
rect 4522 15552 4528 15564
rect 3927 15524 4528 15552
rect 3927 15521 3939 15524
rect 3881 15515 3939 15521
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 6178 15552 6184 15564
rect 5859 15524 6184 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 9048 15552 9076 15648
rect 11514 15580 11520 15632
rect 11572 15620 11578 15632
rect 11790 15620 11796 15632
rect 11572 15592 11796 15620
rect 11572 15580 11578 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 9048 15524 9444 15552
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 4028 15456 4169 15484
rect 4028 15444 4034 15456
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4304 15456 4629 15484
rect 4304 15444 4310 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 5534 15444 5540 15496
rect 5592 15444 5598 15496
rect 8294 15444 8300 15496
rect 8352 15444 8358 15496
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 8536 15456 8677 15484
rect 8536 15444 8542 15456
rect 8665 15453 8677 15456
rect 8711 15453 8723 15487
rect 8665 15447 8723 15453
rect 1762 15376 1768 15428
rect 1820 15376 1826 15428
rect 4065 15419 4123 15425
rect 4065 15385 4077 15419
rect 4111 15416 4123 15419
rect 4706 15416 4712 15428
rect 4111 15388 4712 15416
rect 4111 15385 4123 15388
rect 4065 15379 4123 15385
rect 4706 15376 4712 15388
rect 4764 15416 4770 15428
rect 5261 15419 5319 15425
rect 5261 15416 5273 15419
rect 4764 15388 5273 15416
rect 4764 15376 4770 15388
rect 5261 15385 5273 15388
rect 5307 15385 5319 15419
rect 8680 15416 8708 15447
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9416 15493 9444 15524
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 10100 15524 10425 15552
rect 10100 15512 10106 15524
rect 10413 15521 10425 15524
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15552 10655 15555
rect 11532 15552 11560 15580
rect 10643 15524 11560 15552
rect 10643 15521 10655 15524
rect 10597 15515 10655 15521
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 9088 15456 9137 15484
rect 9088 15444 9094 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 10226 15416 10232 15428
rect 5261 15379 5319 15385
rect 5460 15388 6578 15416
rect 8680 15388 10232 15416
rect 5460 15360 5488 15388
rect 1486 15308 1492 15360
rect 1544 15308 1550 15360
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 4525 15351 4583 15357
rect 4525 15348 4537 15351
rect 4488 15320 4537 15348
rect 4488 15308 4494 15320
rect 4525 15317 4537 15320
rect 4571 15317 4583 15351
rect 4525 15311 4583 15317
rect 5442 15308 5448 15360
rect 5500 15308 5506 15360
rect 5718 15308 5724 15360
rect 5776 15308 5782 15360
rect 6472 15348 6500 15388
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 11164 15416 11192 15447
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11572 15456 11805 15484
rect 11572 15444 11578 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 14642 15444 14648 15496
rect 14700 15444 14706 15496
rect 11164 15388 11836 15416
rect 11808 15360 11836 15388
rect 12066 15376 12072 15428
rect 12124 15376 12130 15428
rect 12526 15376 12532 15428
rect 12584 15376 12590 15428
rect 7098 15348 7104 15360
rect 6472 15320 7104 15348
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 7650 15308 7656 15360
rect 7708 15308 7714 15360
rect 8938 15308 8944 15360
rect 8996 15308 9002 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15348 10011 15351
rect 10318 15348 10324 15360
rect 9999 15320 10324 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 10689 15351 10747 15357
rect 10689 15317 10701 15351
rect 10735 15348 10747 15351
rect 10778 15348 10784 15360
rect 10735 15320 10784 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 11020 15320 11069 15348
rect 11020 15308 11026 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11422 15348 11428 15360
rect 11379 15320 11428 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 11790 15308 11796 15360
rect 11848 15308 11854 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13998 15348 14004 15360
rect 13587 15320 14004 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 14090 15308 14096 15360
rect 14148 15308 14154 15360
rect 1104 15258 16284 15280
rect 1104 15206 3507 15258
rect 3559 15206 3571 15258
rect 3623 15206 3635 15258
rect 3687 15206 3699 15258
rect 3751 15206 3763 15258
rect 3815 15206 7302 15258
rect 7354 15206 7366 15258
rect 7418 15206 7430 15258
rect 7482 15206 7494 15258
rect 7546 15206 7558 15258
rect 7610 15206 11097 15258
rect 11149 15206 11161 15258
rect 11213 15206 11225 15258
rect 11277 15206 11289 15258
rect 11341 15206 11353 15258
rect 11405 15206 14892 15258
rect 14944 15206 14956 15258
rect 15008 15206 15020 15258
rect 15072 15206 15084 15258
rect 15136 15206 15148 15258
rect 15200 15206 16284 15258
rect 1104 15184 16284 15206
rect 4338 15104 4344 15156
rect 4396 15104 4402 15156
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 5258 15144 5264 15156
rect 4479 15116 5264 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 7285 15147 7343 15153
rect 5776 15116 5948 15144
rect 5776 15104 5782 15116
rect 5442 15036 5448 15088
rect 5500 15036 5506 15088
rect 5920 15085 5948 15116
rect 7285 15113 7297 15147
rect 7331 15144 7343 15147
rect 7650 15144 7656 15156
rect 7331 15116 7656 15144
rect 7331 15113 7343 15116
rect 7285 15107 7343 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8938 15144 8944 15156
rect 8036 15116 8944 15144
rect 8036 15085 8064 15116
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 9766 15144 9772 15156
rect 9539 15116 9772 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 11333 15147 11391 15153
rect 10244 15116 11192 15144
rect 5905 15079 5963 15085
rect 5905 15045 5917 15079
rect 5951 15045 5963 15079
rect 8021 15079 8079 15085
rect 5905 15039 5963 15045
rect 6196 15048 7788 15076
rect 6196 15020 6224 15048
rect 3970 14968 3976 15020
rect 4028 14968 4034 15020
rect 6178 14968 6184 15020
rect 6236 14968 6242 15020
rect 7760 15017 7788 15048
rect 8021 15045 8033 15079
rect 8067 15045 8079 15079
rect 9950 15076 9956 15088
rect 9246 15048 9956 15076
rect 8021 15039 8079 15045
rect 9950 15036 9956 15048
rect 10008 15076 10014 15088
rect 10244 15076 10272 15116
rect 11164 15076 11192 15116
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11606 15144 11612 15156
rect 11379 15116 11612 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12526 15144 12532 15156
rect 11716 15116 11928 15144
rect 11716 15076 11744 15116
rect 10008 15048 10350 15076
rect 11164 15048 11744 15076
rect 11900 15076 11928 15116
rect 12176 15116 12532 15144
rect 12176 15076 12204 15116
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15113 13323 15147
rect 13265 15107 13323 15113
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15144 13783 15147
rect 14090 15144 14096 15156
rect 13771 15116 14096 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 13280 15076 13308 15107
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14642 15104 14648 15156
rect 14700 15104 14706 15156
rect 13814 15076 13820 15088
rect 11900 15048 12282 15076
rect 13280 15048 13820 15076
rect 10008 15036 10014 15048
rect 13814 15036 13820 15048
rect 13872 15076 13878 15088
rect 14660 15076 14688 15104
rect 13872 15048 14688 15076
rect 13872 15036 13878 15048
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7193 15011 7251 15017
rect 6779 14980 6868 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14940 2651 14943
rect 2869 14943 2927 14949
rect 2639 14912 2728 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 2700 14816 2728 14912
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 3878 14940 3884 14952
rect 2915 14912 3884 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 6840 14881 6868 14980
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7745 15011 7803 15017
rect 7239 14980 7696 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7377 14943 7435 14949
rect 7377 14940 7389 14943
rect 7064 14912 7389 14940
rect 7064 14900 7070 14912
rect 7377 14909 7389 14912
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 6825 14875 6883 14881
rect 6825 14841 6837 14875
rect 6871 14841 6883 14875
rect 6825 14835 6883 14841
rect 2682 14764 2688 14816
rect 2740 14764 2746 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 7668 14804 7696 14980
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 13136 14980 13952 15008
rect 13136 14968 13142 14980
rect 9585 14943 9643 14949
rect 9585 14940 9597 14943
rect 9324 14912 9597 14940
rect 9324 14816 9352 14912
rect 9585 14909 9597 14912
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 8478 14804 8484 14816
rect 7668 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9306 14764 9312 14816
rect 9364 14764 9370 14816
rect 9600 14804 9628 14903
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 11514 14940 11520 14952
rect 11256 14912 11520 14940
rect 11256 14804 11284 14912
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 13924 14949 13952 14980
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 14056 14980 14749 15008
rect 14056 14968 14062 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11624 14912 11805 14940
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 11624 14872 11652 14912
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 11793 14903 11851 14909
rect 12820 14912 13829 14940
rect 11480 14844 11652 14872
rect 11480 14832 11486 14844
rect 12820 14816 12848 14912
rect 13817 14909 13829 14912
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 13832 14872 13860 14903
rect 14185 14875 14243 14881
rect 14185 14872 14197 14875
rect 13832 14844 14197 14872
rect 14185 14841 14197 14844
rect 14231 14841 14243 14875
rect 14185 14835 14243 14841
rect 9600 14776 11284 14804
rect 12802 14764 12808 14816
rect 12860 14764 12866 14816
rect 13354 14764 13360 14816
rect 13412 14764 13418 14816
rect 1104 14714 16284 14736
rect 1104 14662 2847 14714
rect 2899 14662 2911 14714
rect 2963 14662 2975 14714
rect 3027 14662 3039 14714
rect 3091 14662 3103 14714
rect 3155 14662 6642 14714
rect 6694 14662 6706 14714
rect 6758 14662 6770 14714
rect 6822 14662 6834 14714
rect 6886 14662 6898 14714
rect 6950 14662 10437 14714
rect 10489 14662 10501 14714
rect 10553 14662 10565 14714
rect 10617 14662 10629 14714
rect 10681 14662 10693 14714
rect 10745 14662 14232 14714
rect 14284 14662 14296 14714
rect 14348 14662 14360 14714
rect 14412 14662 14424 14714
rect 14476 14662 14488 14714
rect 14540 14662 16284 14714
rect 1104 14640 16284 14662
rect 3878 14560 3884 14612
rect 3936 14560 3942 14612
rect 4246 14560 4252 14612
rect 4304 14560 4310 14612
rect 5353 14603 5411 14609
rect 5353 14569 5365 14603
rect 5399 14600 5411 14603
rect 5534 14600 5540 14612
rect 5399 14572 5540 14600
rect 5399 14569 5411 14572
rect 5353 14563 5411 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 7006 14600 7012 14612
rect 5644 14572 7012 14600
rect 3605 14535 3663 14541
rect 3605 14501 3617 14535
rect 3651 14532 3663 14535
rect 4264 14532 4292 14560
rect 3651 14504 4292 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 2774 14464 2780 14476
rect 1903 14436 2780 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 5644 14464 5672 14572
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7929 14603 7987 14609
rect 7929 14569 7941 14603
rect 7975 14600 7987 14603
rect 8294 14600 8300 14612
rect 7975 14572 8300 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 9916 14572 10793 14600
rect 9916 14560 9922 14572
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 13814 14600 13820 14612
rect 10781 14563 10839 14569
rect 11440 14572 13820 14600
rect 10318 14492 10324 14544
rect 10376 14532 10382 14544
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 10376 14504 10701 14532
rect 10376 14492 10382 14504
rect 10689 14501 10701 14504
rect 10735 14501 10747 14535
rect 10689 14495 10747 14501
rect 5905 14467 5963 14473
rect 5905 14464 5917 14467
rect 4580 14436 5917 14464
rect 4580 14424 4586 14436
rect 5905 14433 5917 14436
rect 5951 14433 5963 14467
rect 5905 14427 5963 14433
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14464 6515 14467
rect 6546 14464 6552 14476
rect 6503 14436 6552 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9306 14464 9312 14476
rect 8987 14436 9312 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 10284 14436 11253 14464
rect 10284 14424 10290 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 3878 14396 3884 14408
rect 3266 14368 3884 14396
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14396 4123 14399
rect 4246 14396 4252 14408
rect 4111 14368 4252 14396
rect 4111 14365 4123 14368
rect 4065 14359 4123 14365
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4430 14396 4436 14408
rect 4387 14368 4436 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4798 14356 4804 14408
rect 4856 14356 4862 14408
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 6178 14396 6184 14408
rect 5868 14368 6184 14396
rect 5868 14356 5874 14368
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14297 2191 14331
rect 4816 14328 4844 14356
rect 2133 14291 2191 14297
rect 3436 14300 4200 14328
rect 4816 14300 5856 14328
rect 2148 14260 2176 14291
rect 3436 14260 3464 14300
rect 4172 14269 4200 14300
rect 2148 14232 3464 14260
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14229 4215 14263
rect 4157 14223 4215 14229
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4396 14232 4721 14260
rect 4396 14220 4402 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 4709 14223 4767 14229
rect 5169 14263 5227 14269
rect 5169 14229 5181 14263
rect 5215 14260 5227 14263
rect 5534 14260 5540 14272
rect 5215 14232 5540 14260
rect 5215 14229 5227 14232
rect 5169 14223 5227 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5718 14220 5724 14272
rect 5776 14220 5782 14272
rect 5828 14269 5856 14300
rect 5902 14288 5908 14340
rect 5960 14328 5966 14340
rect 5960 14300 6946 14328
rect 5960 14288 5966 14300
rect 9214 14288 9220 14340
rect 9272 14288 9278 14340
rect 9950 14288 9956 14340
rect 10008 14288 10014 14340
rect 11440 14269 11468 14572
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 11532 14436 13921 14464
rect 11532 14408 11560 14436
rect 13909 14433 13921 14436
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 11514 14356 11520 14408
rect 11572 14356 11578 14408
rect 11882 14356 11888 14408
rect 11940 14356 11946 14408
rect 12526 14356 12532 14408
rect 12584 14356 12590 14408
rect 11900 14328 11928 14356
rect 11532 14300 11928 14328
rect 11532 14269 11560 14300
rect 13630 14288 13636 14340
rect 13688 14288 13694 14340
rect 5813 14263 5871 14269
rect 5813 14229 5825 14263
rect 5859 14229 5871 14263
rect 5813 14223 5871 14229
rect 11425 14263 11483 14269
rect 11425 14229 11437 14263
rect 11471 14229 11483 14263
rect 11425 14223 11483 14229
rect 11517 14263 11575 14269
rect 11517 14229 11529 14263
rect 11563 14229 11575 14263
rect 11517 14223 11575 14229
rect 11882 14220 11888 14272
rect 11940 14220 11946 14272
rect 12158 14220 12164 14272
rect 12216 14220 12222 14272
rect 1104 14170 16284 14192
rect 1104 14118 3507 14170
rect 3559 14118 3571 14170
rect 3623 14118 3635 14170
rect 3687 14118 3699 14170
rect 3751 14118 3763 14170
rect 3815 14118 7302 14170
rect 7354 14118 7366 14170
rect 7418 14118 7430 14170
rect 7482 14118 7494 14170
rect 7546 14118 7558 14170
rect 7610 14118 11097 14170
rect 11149 14118 11161 14170
rect 11213 14118 11225 14170
rect 11277 14118 11289 14170
rect 11341 14118 11353 14170
rect 11405 14118 14892 14170
rect 14944 14118 14956 14170
rect 15008 14118 15020 14170
rect 15072 14118 15084 14170
rect 15136 14118 15148 14170
rect 15200 14118 16284 14170
rect 1104 14096 16284 14118
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14025 4307 14059
rect 4249 14019 4307 14025
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 2777 13991 2835 13997
rect 2777 13988 2789 13991
rect 2740 13960 2789 13988
rect 2740 13948 2746 13960
rect 2777 13957 2789 13960
rect 2823 13957 2835 13991
rect 4264 13988 4292 14019
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 5718 14016 5724 14068
rect 5776 14056 5782 14068
rect 5776 14028 6408 14056
rect 5776 14016 5782 14028
rect 6380 14000 6408 14028
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6512 14028 6561 14056
rect 6512 14016 6518 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14056 6975 14059
rect 7650 14056 7656 14068
rect 6963 14028 7656 14056
rect 6963 14025 6975 14028
rect 6917 14019 6975 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9088 14028 9229 14056
rect 9088 14016 9094 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 9766 14056 9772 14068
rect 9723 14028 9772 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 10778 14056 10784 14068
rect 10735 14028 10784 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11790 14056 11796 14068
rect 11563 14028 11796 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 13173 14059 13231 14065
rect 12216 14028 13124 14056
rect 12216 14016 12222 14028
rect 4264 13960 5764 13988
rect 2777 13951 2835 13957
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 5736 13929 5764 13960
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 6420 13960 7021 13988
rect 6420 13948 6426 13960
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 7009 13951 7067 13957
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4856 13892 5181 13920
rect 4856 13880 4862 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 8536 13892 9597 13920
rect 8536 13880 8542 13892
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 11241 13923 11299 13929
rect 11241 13920 11253 13923
rect 10376 13892 11253 13920
rect 10376 13880 10382 13892
rect 11241 13889 11253 13892
rect 11287 13889 11299 13923
rect 11900 13920 11928 14016
rect 12710 13948 12716 14000
rect 12768 13948 12774 14000
rect 12802 13948 12808 14000
rect 12860 13948 12866 14000
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11900 13892 12081 13920
rect 11241 13883 11299 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12636 13892 13032 13920
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2547 13824 2636 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2608 13716 2636 13824
rect 3896 13784 3924 13880
rect 12636 13864 12664 13892
rect 13004 13864 13032 13892
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5074 13852 5080 13864
rect 5031 13824 5080 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5074 13812 5080 13824
rect 5132 13852 5138 13864
rect 7006 13852 7012 13864
rect 5132 13824 7012 13852
rect 5132 13812 5138 13824
rect 7006 13812 7012 13824
rect 7064 13852 7070 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 7064 13824 7113 13852
rect 7064 13812 7070 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 5902 13784 5908 13796
rect 3896 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 9784 13784 9812 13815
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12986 13812 12992 13864
rect 13044 13812 13050 13864
rect 13096 13852 13124 14028
rect 13173 14025 13185 14059
rect 13219 14025 13231 14059
rect 13173 14019 13231 14025
rect 13188 13920 13216 14019
rect 13630 14016 13636 14068
rect 13688 14056 13694 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13688 14028 14013 14056
rect 13688 14016 13694 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14001 14019 14059 14025
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13188 13892 14197 13920
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13096 13824 13829 13852
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 9858 13784 9864 13796
rect 9784 13756 9864 13784
rect 9858 13744 9864 13756
rect 9916 13784 9922 13796
rect 10042 13784 10048 13796
rect 9916 13756 10048 13784
rect 9916 13744 9922 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13265 13787 13323 13793
rect 13265 13784 13277 13787
rect 12860 13756 13277 13784
rect 12860 13744 12866 13756
rect 13265 13753 13277 13756
rect 13311 13753 13323 13787
rect 13265 13747 13323 13753
rect 2774 13716 2780 13728
rect 2608 13688 2780 13716
rect 2774 13676 2780 13688
rect 2832 13716 2838 13728
rect 3234 13716 3240 13728
rect 2832 13688 3240 13716
rect 2832 13676 2838 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4338 13676 4344 13728
rect 4396 13676 4402 13728
rect 1104 13626 16284 13648
rect 1104 13574 2847 13626
rect 2899 13574 2911 13626
rect 2963 13574 2975 13626
rect 3027 13574 3039 13626
rect 3091 13574 3103 13626
rect 3155 13574 6642 13626
rect 6694 13574 6706 13626
rect 6758 13574 6770 13626
rect 6822 13574 6834 13626
rect 6886 13574 6898 13626
rect 6950 13574 10437 13626
rect 10489 13574 10501 13626
rect 10553 13574 10565 13626
rect 10617 13574 10629 13626
rect 10681 13574 10693 13626
rect 10745 13574 14232 13626
rect 14284 13574 14296 13626
rect 14348 13574 14360 13626
rect 14412 13574 14424 13626
rect 14476 13574 14488 13626
rect 14540 13574 16284 13626
rect 1104 13552 16284 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 5074 13472 5080 13524
rect 5132 13472 5138 13524
rect 11793 13515 11851 13521
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 12066 13512 12072 13524
rect 11839 13484 12072 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 13354 13512 13360 13524
rect 12176 13484 13360 13512
rect 5092 13385 5120 13472
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5592 13348 5825 13376
rect 5592 13336 5598 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 12176 13376 12204 13484
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 12897 13447 12955 13453
rect 12897 13413 12909 13447
rect 12943 13413 12955 13447
rect 12897 13407 12955 13413
rect 5813 13339 5871 13345
rect 11624 13348 12204 13376
rect 12345 13379 12403 13385
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 4338 13308 4344 13320
rect 3283 13280 4344 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4798 13268 4804 13320
rect 4856 13268 4862 13320
rect 6546 13268 6552 13320
rect 6604 13268 6610 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 11624 13317 11652 13348
rect 12345 13345 12357 13379
rect 12391 13376 12403 13379
rect 12618 13376 12624 13388
rect 12391 13348 12624 13376
rect 12391 13345 12403 13348
rect 12345 13339 12403 13345
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 12912 13376 12940 13407
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 12912 13348 13553 13376
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 6696 13280 7297 13308
rect 6696 13268 6702 13280
rect 7285 13277 7297 13280
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12115 13280 13001 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 4246 13200 4252 13252
rect 4304 13240 4310 13252
rect 4893 13243 4951 13249
rect 4304 13212 4844 13240
rect 4304 13200 4310 13212
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13172 4491 13175
rect 4706 13172 4712 13184
rect 4479 13144 4712 13172
rect 4479 13141 4491 13144
rect 4433 13135 4491 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4816 13172 4844 13212
rect 4893 13209 4905 13243
rect 4939 13240 4951 13243
rect 6656 13240 6684 13268
rect 4939 13212 6684 13240
rect 12529 13243 12587 13249
rect 4939 13209 4951 13212
rect 4893 13203 4951 13209
rect 12529 13209 12541 13243
rect 12575 13240 12587 13243
rect 12710 13240 12716 13252
rect 12575 13212 12716 13240
rect 12575 13209 12587 13212
rect 12529 13203 12587 13209
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 4816 13144 5273 13172
rect 5261 13141 5273 13144
rect 5307 13141 5319 13175
rect 5261 13135 5319 13141
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5776 13144 6009 13172
rect 5776 13132 5782 13144
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 6730 13132 6736 13184
rect 6788 13132 6794 13184
rect 11882 13132 11888 13184
rect 11940 13132 11946 13184
rect 12434 13132 12440 13184
rect 12492 13132 12498 13184
rect 1104 13082 16284 13104
rect 1104 13030 3507 13082
rect 3559 13030 3571 13082
rect 3623 13030 3635 13082
rect 3687 13030 3699 13082
rect 3751 13030 3763 13082
rect 3815 13030 7302 13082
rect 7354 13030 7366 13082
rect 7418 13030 7430 13082
rect 7482 13030 7494 13082
rect 7546 13030 7558 13082
rect 7610 13030 11097 13082
rect 11149 13030 11161 13082
rect 11213 13030 11225 13082
rect 11277 13030 11289 13082
rect 11341 13030 11353 13082
rect 11405 13030 14892 13082
rect 14944 13030 14956 13082
rect 15008 13030 15020 13082
rect 15072 13030 15084 13082
rect 15136 13030 15148 13082
rect 15200 13030 16284 13082
rect 1104 13008 16284 13030
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 6365 12971 6423 12977
rect 6365 12937 6377 12971
rect 6411 12968 6423 12971
rect 6546 12968 6552 12980
rect 6411 12940 6552 12968
rect 6411 12937 6423 12940
rect 6365 12931 6423 12937
rect 5828 12900 5856 12931
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 6638 12928 6644 12980
rect 6696 12928 6702 12980
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 12492 12940 13277 12968
rect 12492 12928 12498 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 6656 12900 6684 12928
rect 5828 12872 6684 12900
rect 11793 12903 11851 12909
rect 11793 12869 11805 12903
rect 11839 12900 11851 12903
rect 11900 12900 11928 12928
rect 11839 12872 11928 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 12526 12860 12532 12912
rect 12584 12860 12590 12912
rect 5902 12832 5908 12844
rect 5474 12804 5908 12832
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7558 12832 7564 12844
rect 6871 12804 7564 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 13280 12832 13308 12931
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13280 12804 13921 12832
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 13909 12795 13967 12801
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3292 12736 4077 12764
rect 3292 12724 3298 12736
rect 4065 12733 4077 12736
rect 4111 12733 4123 12767
rect 4065 12727 4123 12733
rect 4338 12724 4344 12776
rect 4396 12724 4402 12776
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7834 12764 7840 12776
rect 7064 12736 7840 12764
rect 7064 12724 7070 12736
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 13354 12588 13360 12640
rect 13412 12588 13418 12640
rect 1104 12538 16284 12560
rect 1104 12486 2847 12538
rect 2899 12486 2911 12538
rect 2963 12486 2975 12538
rect 3027 12486 3039 12538
rect 3091 12486 3103 12538
rect 3155 12486 6642 12538
rect 6694 12486 6706 12538
rect 6758 12486 6770 12538
rect 6822 12486 6834 12538
rect 6886 12486 6898 12538
rect 6950 12486 10437 12538
rect 10489 12486 10501 12538
rect 10553 12486 10565 12538
rect 10617 12486 10629 12538
rect 10681 12486 10693 12538
rect 10745 12486 14232 12538
rect 14284 12486 14296 12538
rect 14348 12486 14360 12538
rect 14412 12486 14424 12538
rect 14476 12486 14488 12538
rect 14540 12486 16284 12538
rect 1104 12464 16284 12486
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4338 12424 4344 12436
rect 4295 12396 4344 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9916 12396 12020 12424
rect 9916 12384 9922 12396
rect 11425 12359 11483 12365
rect 11425 12325 11437 12359
rect 11471 12325 11483 12359
rect 11425 12319 11483 12325
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 2225 12291 2283 12297
rect 2225 12288 2237 12291
rect 1820 12260 2237 12288
rect 1820 12248 1826 12260
rect 2225 12257 2237 12260
rect 2271 12257 2283 12291
rect 2225 12251 2283 12257
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4764 12260 5089 12288
rect 4764 12248 4770 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 6086 12288 6092 12300
rect 5868 12260 6092 12288
rect 5868 12248 5874 12260
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 7558 12248 7564 12300
rect 7616 12288 7622 12300
rect 8018 12288 8024 12300
rect 7616 12260 8024 12288
rect 7616 12248 7622 12260
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11440 12288 11468 12319
rect 11992 12297 12020 12396
rect 11379 12260 11468 12288
rect 11977 12291 12035 12297
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12618 12288 12624 12300
rect 12023 12260 12624 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3326 12220 3332 12232
rect 3191 12192 3332 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4479 12192 4537 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9732 12192 9781 12220
rect 9732 12180 9738 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 13354 12220 13360 12232
rect 11839 12192 13360 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 14642 12180 14648 12232
rect 14700 12180 14706 12232
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14792 12192 15025 12220
rect 14792 12180 14798 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15838 12180 15844 12232
rect 15896 12180 15902 12232
rect 6089 12155 6147 12161
rect 6089 12152 6101 12155
rect 5736 12124 6101 12152
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 2869 12087 2927 12093
rect 2869 12084 2881 12087
rect 2740 12056 2881 12084
rect 2740 12044 2746 12056
rect 2869 12053 2881 12056
rect 2915 12053 2927 12087
rect 2869 12047 2927 12053
rect 2958 12044 2964 12096
rect 3016 12044 3022 12096
rect 5736 12093 5764 12124
rect 6089 12121 6101 12124
rect 6135 12121 6147 12155
rect 6089 12115 6147 12121
rect 5721 12087 5779 12093
rect 5721 12053 5733 12087
rect 5767 12053 5779 12087
rect 5721 12047 5779 12053
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7208 12084 7236 12180
rect 7064 12056 7236 12084
rect 7064 12044 7070 12056
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7432 12056 7665 12084
rect 7432 12044 7438 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8444 12056 9229 12084
rect 8444 12044 8450 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11885 12087 11943 12093
rect 11885 12084 11897 12087
rect 11848 12056 11897 12084
rect 11848 12044 11854 12056
rect 11885 12053 11897 12056
rect 11931 12053 11943 12087
rect 11885 12047 11943 12053
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13596 12056 14105 12084
rect 13596 12044 13602 12056
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 14550 12044 14556 12096
rect 14608 12084 14614 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14608 12056 14841 12084
rect 14608 12044 14614 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 14829 12047 14887 12053
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 1104 11994 16284 12016
rect 1104 11942 3507 11994
rect 3559 11942 3571 11994
rect 3623 11942 3635 11994
rect 3687 11942 3699 11994
rect 3751 11942 3763 11994
rect 3815 11942 7302 11994
rect 7354 11942 7366 11994
rect 7418 11942 7430 11994
rect 7482 11942 7494 11994
rect 7546 11942 7558 11994
rect 7610 11942 11097 11994
rect 11149 11942 11161 11994
rect 11213 11942 11225 11994
rect 11277 11942 11289 11994
rect 11341 11942 11353 11994
rect 11405 11942 14892 11994
rect 14944 11942 14956 11994
rect 15008 11942 15020 11994
rect 15072 11942 15084 11994
rect 15136 11942 15148 11994
rect 15200 11942 16284 11994
rect 1104 11920 16284 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 1670 11880 1676 11892
rect 1535 11852 1676 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 2530 11784 3464 11812
rect 3436 11756 3464 11784
rect 3418 11704 3424 11756
rect 3476 11704 3482 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 6932 11744 6960 11843
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 7248 11852 7297 11880
rect 7248 11840 7254 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 7377 11883 7435 11889
rect 7377 11849 7389 11883
rect 7423 11880 7435 11883
rect 7423 11852 7696 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 6687 11716 6960 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7668 11744 7696 11852
rect 10686 11840 10692 11892
rect 10744 11840 10750 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 12851 11852 13216 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 8478 11812 8484 11824
rect 8312 11784 8484 11812
rect 8312 11744 8340 11784
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 10505 11815 10563 11821
rect 10505 11812 10517 11815
rect 9916 11784 10517 11812
rect 9916 11772 9922 11784
rect 10505 11781 10517 11784
rect 10551 11781 10563 11815
rect 10505 11775 10563 11781
rect 9950 11744 9956 11756
rect 7248 11716 7512 11744
rect 7668 11716 8340 11744
rect 9706 11716 9956 11744
rect 7248 11704 7254 11716
rect 2958 11636 2964 11688
rect 3016 11636 3022 11688
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 7484 11685 7512 11716
rect 9950 11704 9956 11716
rect 10008 11744 10014 11756
rect 10704 11744 10732 11840
rect 13188 11821 13216 11852
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 14734 11840 14740 11892
rect 14792 11840 14798 11892
rect 13173 11815 13231 11821
rect 13173 11781 13185 11815
rect 13219 11781 13231 11815
rect 15286 11812 15292 11824
rect 13173 11775 13231 11781
rect 15212 11784 15292 11812
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10008 11716 10272 11744
rect 10704 11716 11253 11744
rect 10008 11704 10014 11716
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 3252 11608 3280 11636
rect 6086 11608 6092 11620
rect 3252 11580 6092 11608
rect 6086 11568 6092 11580
rect 6144 11608 6150 11620
rect 8312 11608 8340 11639
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 6144 11580 8340 11608
rect 6144 11568 6150 11580
rect 6454 11500 6460 11552
rect 6512 11500 6518 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 10244 11549 10272 11716
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 14734 11744 14740 11756
rect 14306 11716 14740 11744
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 12342 11676 12348 11688
rect 11572 11648 12348 11676
rect 11572 11636 11578 11648
rect 12342 11636 12348 11648
rect 12400 11676 12406 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12400 11648 12909 11676
rect 12400 11636 12406 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13538 11636 13544 11688
rect 13596 11676 13602 11688
rect 15120 11676 15148 11707
rect 15212 11685 15240 11784
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 13596 11648 15148 11676
rect 15197 11679 15255 11685
rect 13596 11636 13602 11648
rect 15197 11645 15209 11679
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 9732 11512 10057 11540
rect 9732 11500 9738 11512
rect 10045 11509 10057 11512
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 10229 11543 10287 11549
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10318 11540 10324 11552
rect 10275 11512 10324 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10928 11512 11069 11540
rect 10928 11500 10934 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 15212 11540 15240 11639
rect 15378 11636 15384 11688
rect 15436 11636 15442 11688
rect 14700 11512 15240 11540
rect 14700 11500 14706 11512
rect 1104 11450 16284 11472
rect 1104 11398 2847 11450
rect 2899 11398 2911 11450
rect 2963 11398 2975 11450
rect 3027 11398 3039 11450
rect 3091 11398 3103 11450
rect 3155 11398 6642 11450
rect 6694 11398 6706 11450
rect 6758 11398 6770 11450
rect 6822 11398 6834 11450
rect 6886 11398 6898 11450
rect 6950 11398 10437 11450
rect 10489 11398 10501 11450
rect 10553 11398 10565 11450
rect 10617 11398 10629 11450
rect 10681 11398 10693 11450
rect 10745 11398 14232 11450
rect 14284 11398 14296 11450
rect 14348 11398 14360 11450
rect 14412 11398 14424 11450
rect 14476 11398 14488 11450
rect 14540 11398 16284 11450
rect 1104 11376 16284 11398
rect 2774 11296 2780 11348
rect 2832 11296 2838 11348
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3326 11336 3332 11348
rect 3283 11308 3332 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 6076 11339 6134 11345
rect 6076 11305 6088 11339
rect 6122 11336 6134 11339
rect 6454 11336 6460 11348
rect 6122 11308 6460 11336
rect 6122 11305 6134 11308
rect 6076 11299 6134 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7742 11336 7748 11348
rect 7607 11308 7748 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7742 11296 7748 11308
rect 7800 11336 7806 11348
rect 8202 11336 8208 11348
rect 7800 11308 8208 11336
rect 7800 11296 7806 11308
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8628 11308 8953 11336
rect 8628 11296 8634 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 10768 11339 10826 11345
rect 10768 11305 10780 11339
rect 10814 11336 10826 11339
rect 10870 11336 10876 11348
rect 10814 11308 10876 11336
rect 10814 11305 10826 11308
rect 10768 11299 10826 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11020 11308 12434 11336
rect 11020 11296 11026 11308
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2700 11064 2728 11163
rect 2792 11132 2820 11296
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 6086 11200 6092 11212
rect 5859 11172 6092 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 8294 11200 8300 11212
rect 8251 11172 8300 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8404 11141 8432 11296
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2792 11104 2881 11132
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8772 11132 8800 11231
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 11514 11200 11520 11212
rect 10551 11172 11520 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11808 11172 12265 11200
rect 11808 11144 11836 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12406 11200 12434 11308
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12676 11308 13093 11336
rect 12676 11296 12682 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 14356 11339 14414 11345
rect 14356 11305 14368 11339
rect 14402 11336 14414 11339
rect 14550 11336 14556 11348
rect 14402 11308 14556 11336
rect 14402 11305 14414 11308
rect 14356 11299 14414 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15838 11296 15844 11348
rect 15896 11296 15902 11348
rect 12989 11271 13047 11277
rect 12989 11237 13001 11271
rect 13035 11268 13047 11271
rect 13814 11268 13820 11280
rect 13035 11240 13820 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 12406 11172 13492 11200
rect 12253 11163 12311 11169
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8772 11104 9137 11132
rect 8389 11095 8447 11101
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 9784 11104 9873 11132
rect 3142 11064 3148 11076
rect 2700 11036 3148 11064
rect 3142 11024 3148 11036
rect 3200 11024 3206 11076
rect 6362 11064 6368 11076
rect 5920 11036 6368 11064
rect 5920 11008 5948 11036
rect 6362 11024 6368 11036
rect 6420 11064 6426 11076
rect 9324 11064 9352 11092
rect 9784 11076 9812 11104
rect 9861 11101 9873 11104
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 11790 11092 11796 11144
rect 11848 11092 11854 11144
rect 12526 11132 12532 11144
rect 11914 11104 12532 11132
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 13464 11141 13492 11172
rect 13538 11160 13544 11212
rect 13596 11160 13602 11212
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 15378 11200 15384 11212
rect 13679 11172 15384 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 6420 11036 6578 11064
rect 8220 11036 9352 11064
rect 6420 11024 6426 11036
rect 8220 11008 8248 11036
rect 9766 11024 9772 11076
rect 9824 11024 9830 11076
rect 12820 11064 12848 11095
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13780 11104 14105 11132
rect 13780 11092 13786 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 13906 11064 13912 11076
rect 10336 11036 11192 11064
rect 12820 11036 13912 11064
rect 2774 10956 2780 11008
rect 2832 10956 2838 11008
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 8202 10956 8208 11008
rect 8260 10956 8266 11008
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8478 10996 8484 11008
rect 8343 10968 8484 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8478 10956 8484 10968
rect 8536 10996 8542 11008
rect 9950 10996 9956 11008
rect 8536 10968 9956 10996
rect 8536 10956 8542 10968
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10336 11005 10364 11036
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10965 10379 10999
rect 11164 10996 11192 11036
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14752 11036 14858 11064
rect 14752 11008 14780 11036
rect 11422 10996 11428 11008
rect 11164 10968 11428 10996
rect 10321 10959 10379 10965
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 1104 10906 16284 10928
rect 1104 10854 3507 10906
rect 3559 10854 3571 10906
rect 3623 10854 3635 10906
rect 3687 10854 3699 10906
rect 3751 10854 3763 10906
rect 3815 10854 7302 10906
rect 7354 10854 7366 10906
rect 7418 10854 7430 10906
rect 7482 10854 7494 10906
rect 7546 10854 7558 10906
rect 7610 10854 11097 10906
rect 11149 10854 11161 10906
rect 11213 10854 11225 10906
rect 11277 10854 11289 10906
rect 11341 10854 11353 10906
rect 11405 10854 14892 10906
rect 14944 10854 14956 10906
rect 15008 10854 15020 10906
rect 15072 10854 15084 10906
rect 15136 10854 15148 10906
rect 15200 10854 16284 10906
rect 1104 10832 16284 10854
rect 3234 10792 3240 10804
rect 2240 10764 3240 10792
rect 2240 10665 2268 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 7190 10752 7196 10804
rect 7248 10752 7254 10804
rect 3510 10684 3516 10736
rect 3568 10684 3574 10736
rect 4525 10727 4583 10733
rect 4525 10693 4537 10727
rect 4571 10724 4583 10727
rect 5902 10724 5908 10736
rect 4571 10696 5908 10724
rect 4571 10693 4583 10696
rect 4525 10687 4583 10693
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2498 10548 2504 10600
rect 2556 10548 2562 10600
rect 3528 10588 3556 10684
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4338 10656 4344 10668
rect 4203 10628 4344 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4540 10588 4568 10687
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 7055 10696 8800 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 8772 10668 8800 10696
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9766 10724 9772 10736
rect 9272 10696 9772 10724
rect 9272 10684 9278 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 10318 10684 10324 10736
rect 10376 10684 10382 10736
rect 11057 10727 11115 10733
rect 11057 10693 11069 10727
rect 11103 10724 11115 10727
rect 11422 10724 11428 10736
rect 11103 10696 11428 10724
rect 11103 10693 11115 10696
rect 11057 10687 11115 10693
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 13722 10724 13728 10736
rect 13556 10696 13728 10724
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 3528 10560 4568 10588
rect 7116 10628 7297 10656
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 6604 10492 6653 10520
rect 6604 10480 6610 10492
rect 6641 10489 6653 10492
rect 6687 10489 6699 10523
rect 6641 10483 6699 10489
rect 7116 10464 7144 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7650 10616 7656 10668
rect 7708 10616 7714 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8202 10656 8208 10668
rect 8067 10628 8208 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 7190 10548 7196 10600
rect 7248 10588 7254 10600
rect 8036 10588 8064 10619
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 7248 10560 8064 10588
rect 8404 10588 8432 10619
rect 8754 10616 8760 10668
rect 8812 10616 8818 10668
rect 9398 10656 9404 10668
rect 8864 10628 9404 10656
rect 8864 10588 8892 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 11333 10659 11391 10665
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 12342 10656 12348 10668
rect 11379 10628 12348 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 12342 10616 12348 10628
rect 12400 10656 12406 10668
rect 13446 10656 13452 10668
rect 12400 10628 13452 10656
rect 12400 10616 12406 10628
rect 13446 10616 13452 10628
rect 13504 10656 13510 10668
rect 13556 10665 13584 10696
rect 13722 10684 13728 10696
rect 13780 10684 13786 10736
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13504 10628 13553 10656
rect 13504 10616 13510 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 14884 10628 14950 10656
rect 14884 10616 14890 10628
rect 8404 10560 8892 10588
rect 8941 10591 8999 10597
rect 7248 10548 7254 10560
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 8987 10560 9628 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 3970 10412 3976 10464
rect 4028 10412 4034 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7098 10452 7104 10464
rect 7055 10424 7104 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 9490 10412 9496 10464
rect 9548 10412 9554 10464
rect 9600 10461 9628 10560
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 10042 10452 10048 10464
rect 9631 10424 10048 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 15286 10412 15292 10464
rect 15344 10412 15350 10464
rect 1104 10362 16284 10384
rect 1104 10310 2847 10362
rect 2899 10310 2911 10362
rect 2963 10310 2975 10362
rect 3027 10310 3039 10362
rect 3091 10310 3103 10362
rect 3155 10310 6642 10362
rect 6694 10310 6706 10362
rect 6758 10310 6770 10362
rect 6822 10310 6834 10362
rect 6886 10310 6898 10362
rect 6950 10310 10437 10362
rect 10489 10310 10501 10362
rect 10553 10310 10565 10362
rect 10617 10310 10629 10362
rect 10681 10310 10693 10362
rect 10745 10310 14232 10362
rect 14284 10310 14296 10362
rect 14348 10310 14360 10362
rect 14412 10310 14424 10362
rect 14476 10310 14488 10362
rect 14540 10310 16284 10362
rect 1104 10288 16284 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10217 2191 10251
rect 2133 10211 2191 10217
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2498 10248 2504 10260
rect 2271 10220 2504 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2148 10180 2176 10211
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 3970 10248 3976 10260
rect 2608 10220 3976 10248
rect 2608 10180 2636 10220
rect 2148 10152 2636 10180
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3513 10115 3571 10121
rect 2731 10084 3464 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2038 10004 2044 10056
rect 2096 10004 2102 10056
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 2314 10044 2320 10056
rect 2179 10016 2320 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2639 10016 2881 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 3436 10044 3464 10084
rect 3513 10081 3525 10115
rect 3559 10112 3571 10115
rect 3620 10112 3648 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 6086 10248 6092 10260
rect 5767 10220 6092 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7742 10208 7748 10260
rect 7800 10208 7806 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8352 10220 8953 10248
rect 8352 10208 8358 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9214 10248 9220 10260
rect 9171 10220 9220 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 8021 10183 8079 10189
rect 8021 10180 8033 10183
rect 3559 10084 3648 10112
rect 3712 10152 8033 10180
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 3712 10044 3740 10152
rect 8021 10149 8033 10152
rect 8067 10149 8079 10183
rect 8021 10143 8079 10149
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9140 10180 9168 10211
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10192 10220 10333 10248
rect 10192 10208 10198 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12342 10248 12348 10260
rect 11931 10220 12348 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13964 10220 14289 10248
rect 13964 10208 13970 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 15378 10208 15384 10260
rect 15436 10208 15442 10260
rect 8536 10152 9168 10180
rect 9508 10180 9536 10208
rect 9508 10152 9904 10180
rect 8536 10140 8542 10152
rect 4522 10072 4528 10124
rect 4580 10072 4586 10124
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 5031 10084 7113 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7742 10112 7748 10124
rect 7101 10075 7159 10081
rect 7392 10084 7748 10112
rect 3436 10016 3740 10044
rect 2869 10007 2927 10013
rect 3878 10004 3884 10056
rect 3936 10004 3942 10056
rect 7392 10053 7420 10084
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8665 10115 8723 10121
rect 8220 10084 8432 10112
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4479 10016 4905 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7650 10044 7656 10056
rect 7515 10016 7656 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8220 10044 8248 10084
rect 7883 10016 8248 10044
rect 8297 10047 8355 10053
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8297 10013 8309 10047
rect 8343 10013 8355 10047
rect 8404 10044 8432 10084
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 9674 10112 9680 10124
rect 8711 10084 9680 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 9876 10121 9904 10152
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 15105 10183 15163 10189
rect 15105 10180 15117 10183
rect 14148 10152 15117 10180
rect 14148 10140 14154 10152
rect 15105 10149 15117 10152
rect 15151 10149 15163 10183
rect 15105 10143 15163 10149
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10081 9919 10115
rect 9861 10075 9919 10081
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 14608 10084 14933 10112
rect 14608 10072 14614 10084
rect 14921 10081 14933 10084
rect 14967 10112 14979 10115
rect 15396 10112 15424 10208
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 14967 10084 15669 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 8404 10016 8769 10044
rect 8297 10007 8355 10013
rect 8757 10013 8769 10016
rect 8803 10044 8815 10047
rect 9214 10044 9220 10056
rect 8803 10016 9220 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 8202 9976 8208 9988
rect 7055 9948 8208 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9908 1823 9911
rect 2774 9908 2780 9920
rect 1811 9880 2780 9908
rect 1811 9877 1823 9880
rect 1765 9871 1823 9877
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7098 9908 7104 9920
rect 6972 9880 7104 9908
rect 6972 9868 6978 9880
rect 7098 9868 7104 9880
rect 7156 9908 7162 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7156 9880 7573 9908
rect 7156 9868 7162 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 8110 9908 8116 9920
rect 7800 9880 8116 9908
rect 7800 9868 7806 9880
rect 8110 9868 8116 9880
rect 8168 9908 8174 9920
rect 8312 9908 8340 10007
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9490 10004 9496 10056
rect 9548 10004 9554 10056
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 10376 10016 10425 10044
rect 10376 10004 10382 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10962 10004 10968 10056
rect 11020 10004 11026 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 8389 9979 8447 9985
rect 8389 9945 8401 9979
rect 8435 9976 8447 9979
rect 10594 9976 10600 9988
rect 8435 9948 10600 9976
rect 8435 9945 8447 9948
rect 8389 9939 8447 9945
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 8168 9880 8340 9908
rect 8168 9868 8174 9880
rect 8478 9868 8484 9920
rect 8536 9868 8542 9920
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 8812 9880 9137 9908
rect 8812 9868 8818 9880
rect 9125 9877 9137 9880
rect 9171 9877 9183 9911
rect 9125 9871 9183 9877
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10980 9908 11008 10004
rect 10008 9880 11008 9908
rect 14737 9911 14795 9917
rect 10008 9868 10014 9880
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 15470 9908 15476 9920
rect 14783 9880 15476 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15562 9868 15568 9920
rect 15620 9868 15626 9920
rect 1104 9818 16284 9840
rect 1104 9766 3507 9818
rect 3559 9766 3571 9818
rect 3623 9766 3635 9818
rect 3687 9766 3699 9818
rect 3751 9766 3763 9818
rect 3815 9766 7302 9818
rect 7354 9766 7366 9818
rect 7418 9766 7430 9818
rect 7482 9766 7494 9818
rect 7546 9766 7558 9818
rect 7610 9766 11097 9818
rect 11149 9766 11161 9818
rect 11213 9766 11225 9818
rect 11277 9766 11289 9818
rect 11341 9766 11353 9818
rect 11405 9766 14892 9818
rect 14944 9766 14956 9818
rect 15008 9766 15020 9818
rect 15072 9766 15084 9818
rect 15136 9766 15148 9818
rect 15200 9766 16284 9818
rect 1104 9744 16284 9766
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 2409 9707 2467 9713
rect 2409 9704 2421 9707
rect 2096 9676 2421 9704
rect 2096 9664 2102 9676
rect 2409 9673 2421 9676
rect 2455 9704 2467 9707
rect 3786 9704 3792 9716
rect 2455 9676 3792 9704
rect 2455 9673 2467 9676
rect 2409 9667 2467 9673
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 7098 9704 7104 9716
rect 4396 9676 7104 9704
rect 4396 9664 4402 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 7469 9707 7527 9713
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7650 9704 7656 9716
rect 7515 9676 7656 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 10318 9704 10324 9716
rect 9600 9676 10324 9704
rect 3418 9596 3424 9648
rect 3476 9596 3482 9648
rect 3881 9639 3939 9645
rect 3881 9605 3893 9639
rect 3927 9636 3939 9639
rect 4522 9636 4528 9648
rect 3927 9608 4528 9636
rect 3927 9605 3939 9608
rect 3881 9599 3939 9605
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 6546 9596 6552 9648
rect 6604 9596 6610 9648
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 7208 9636 7236 9664
rect 6779 9608 7236 9636
rect 7668 9608 8248 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6564 9568 6592 9596
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6135 9540 6408 9568
rect 6564 9540 6837 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4522 9500 4528 9512
rect 4203 9472 4528 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4939 9472 4997 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 4985 9469 4997 9472
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5442 9460 5448 9512
rect 5500 9460 5506 9512
rect 6380 9441 6408 9540
rect 6825 9537 6837 9540
rect 6871 9568 6883 9571
rect 7190 9568 7196 9580
rect 6871 9540 7196 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7668 9577 7696 9608
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 6365 9435 6423 9441
rect 6365 9401 6377 9435
rect 6411 9401 6423 9435
rect 6365 9395 6423 9401
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 3752 9336 4261 9364
rect 3752 9324 3758 9336
rect 4249 9333 4261 9336
rect 4295 9333 4307 9367
rect 4249 9327 4307 9333
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5868 9336 5917 9364
rect 5868 9324 5874 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 7024 9364 7052 9463
rect 7760 9432 7788 9531
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 8220 9568 8248 9608
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8352 9608 8953 9636
rect 8352 9596 8358 9608
rect 8941 9605 8953 9608
rect 8987 9636 8999 9639
rect 9600 9636 9628 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10594 9664 10600 9716
rect 10652 9664 10658 9716
rect 14090 9664 14096 9716
rect 14148 9664 14154 9716
rect 15470 9664 15476 9716
rect 15528 9704 15534 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15528 9676 15945 9704
rect 15528 9664 15534 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 14108 9636 14136 9664
rect 8987 9608 9628 9636
rect 13188 9608 14136 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 8386 9568 8392 9580
rect 8220 9540 8392 9568
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 8570 9568 8576 9580
rect 8527 9540 8576 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9490 9568 9496 9580
rect 8720 9540 9496 9568
rect 8720 9528 8726 9540
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8202 9500 8208 9512
rect 7975 9472 8208 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8202 9460 8208 9472
rect 8260 9500 8266 9512
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 8260 9472 8309 9500
rect 8260 9460 8266 9472
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 8404 9500 8432 9528
rect 10134 9500 10140 9512
rect 8404 9472 10140 9500
rect 8297 9463 8355 9469
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 10796 9500 10824 9531
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11790 9568 11796 9580
rect 11195 9540 11796 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 13188 9577 13216 9608
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 10192 9472 10824 9500
rect 10192 9460 10198 9472
rect 13446 9460 13452 9512
rect 13504 9460 13510 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13556 9472 13737 9500
rect 8478 9432 8484 9444
rect 7760 9404 8484 9432
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 13357 9435 13415 9441
rect 13357 9401 13369 9435
rect 13403 9432 13415 9435
rect 13556 9432 13584 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14734 9500 14740 9512
rect 13872 9472 14740 9500
rect 13872 9460 13878 9472
rect 14734 9460 14740 9472
rect 14792 9500 14798 9512
rect 14844 9500 14872 9554
rect 15286 9528 15292 9580
rect 15344 9528 15350 9580
rect 14792 9472 14872 9500
rect 14792 9460 14798 9472
rect 13403 9404 13584 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 6604 9336 7052 9364
rect 6604 9324 6610 9336
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 10962 9364 10968 9376
rect 8168 9336 10968 9364
rect 8168 9324 8174 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11238 9364 11244 9376
rect 11103 9336 11244 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15286 9364 15292 9376
rect 15243 9336 15292 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 1104 9274 16284 9296
rect 1104 9222 2847 9274
rect 2899 9222 2911 9274
rect 2963 9222 2975 9274
rect 3027 9222 3039 9274
rect 3091 9222 3103 9274
rect 3155 9222 6642 9274
rect 6694 9222 6706 9274
rect 6758 9222 6770 9274
rect 6822 9222 6834 9274
rect 6886 9222 6898 9274
rect 6950 9222 10437 9274
rect 10489 9222 10501 9274
rect 10553 9222 10565 9274
rect 10617 9222 10629 9274
rect 10681 9222 10693 9274
rect 10745 9222 14232 9274
rect 14284 9222 14296 9274
rect 14348 9222 14360 9274
rect 14412 9222 14424 9274
rect 14476 9222 14488 9274
rect 14540 9222 16284 9274
rect 1104 9200 16284 9222
rect 1857 9163 1915 9169
rect 1857 9129 1869 9163
rect 1903 9160 1915 9163
rect 2314 9160 2320 9172
rect 1903 9132 2320 9160
rect 1903 9129 1915 9132
rect 1857 9123 1915 9129
rect 2314 9120 2320 9132
rect 2372 9160 2378 9172
rect 4433 9163 4491 9169
rect 2372 9132 3832 9160
rect 2372 9120 2378 9132
rect 3694 9052 3700 9104
rect 3752 9052 3758 9104
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3712 9024 3740 9052
rect 3804 9033 3832 9132
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 5350 9160 5356 9172
rect 4479 9132 5356 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 8220 9132 8309 9160
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 7377 9095 7435 9101
rect 7377 9092 7389 9095
rect 6880 9064 7389 9092
rect 6880 9052 6886 9064
rect 7377 9061 7389 9064
rect 7423 9061 7435 9095
rect 7377 9055 7435 9061
rect 3375 8996 3740 9024
rect 3789 9027 3847 9033
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3789 8993 3801 9027
rect 3835 8993 3847 9027
rect 3789 8987 3847 8993
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 5810 9024 5816 9036
rect 5767 8996 5816 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 6788 8996 7941 9024
rect 6788 8984 6794 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 8220 9024 8248 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8444 9132 8677 9160
rect 8444 9120 8450 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 9272 9132 9505 9160
rect 9272 9120 9278 9132
rect 8570 9024 8576 9036
rect 7929 8987 7987 8993
rect 8128 8996 8576 9024
rect 8128 8968 8156 8996
rect 8570 8984 8576 8996
rect 8628 9024 8634 9036
rect 9309 9027 9367 9033
rect 8628 8996 9260 9024
rect 8628 8984 8634 8996
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 3605 8919 3663 8925
rect 4540 8928 5457 8956
rect 3326 8888 3332 8900
rect 2898 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 3620 8820 3648 8919
rect 4540 8832 4568 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 7190 8916 7196 8968
rect 7248 8916 7254 8968
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8110 8956 8116 8968
rect 7883 8928 8116 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8662 8956 8668 8968
rect 8251 8928 8668 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 6454 8848 6460 8900
rect 6512 8848 6518 8900
rect 4522 8820 4528 8832
rect 3620 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 7208 8829 7236 8916
rect 7742 8848 7748 8900
rect 7800 8848 7806 8900
rect 7193 8823 7251 8829
rect 7193 8789 7205 8823
rect 7239 8820 7251 8823
rect 8312 8820 8340 8928
rect 8662 8916 8668 8928
rect 8720 8956 8726 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8720 8928 9137 8956
rect 8720 8916 8726 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9232 8956 9260 8996
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 9416 9024 9444 9132
rect 9493 9129 9505 9132
rect 9539 9129 9551 9163
rect 9493 9123 9551 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9824 9132 10609 9160
rect 9824 9120 9830 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9129 10839 9163
rect 10781 9123 10839 9129
rect 10796 9092 10824 9123
rect 14550 9120 14556 9172
rect 14608 9120 14614 9172
rect 9784 9064 10824 9092
rect 12529 9095 12587 9101
rect 9355 8996 9536 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 9232 8928 9413 8956
rect 9125 8919 9183 8925
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 7239 8792 8340 8820
rect 8941 8823 8999 8829
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 8941 8789 8953 8823
rect 8987 8820 8999 8823
rect 9214 8820 9220 8832
rect 8987 8792 9220 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9508 8820 9536 8996
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 9784 9024 9812 9064
rect 12529 9061 12541 9095
rect 12575 9092 12587 9095
rect 14568 9092 14596 9120
rect 12575 9064 14596 9092
rect 14829 9095 14887 9101
rect 12575 9061 12587 9064
rect 12529 9055 12587 9061
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 9732 8996 9812 9024
rect 9968 8996 10885 9024
rect 9732 8984 9738 8996
rect 9600 8888 9628 8984
rect 9968 8965 9996 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 14292 9033 14320 9064
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 15378 9092 15384 9104
rect 14875 9064 15384 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 14240 8996 14289 9024
rect 14240 8984 14246 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 15654 9024 15660 9036
rect 14277 8987 14335 8993
rect 14476 8996 15660 9024
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9784 8928 9965 8956
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 9600 8860 9689 8888
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 9677 8851 9735 8857
rect 9784 8820 9812 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10152 8888 10180 8919
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10284 8928 10333 8956
rect 10284 8916 10290 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10744 8928 10977 8956
rect 10744 8916 10750 8928
rect 10965 8925 10977 8928
rect 11011 8956 11023 8959
rect 11057 8959 11115 8965
rect 11057 8956 11069 8959
rect 11011 8928 11069 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11057 8925 11069 8928
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 11471 8928 12357 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 14476 8965 14504 8996
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 15470 8916 15476 8968
rect 15528 8916 15534 8968
rect 10778 8888 10784 8900
rect 10152 8860 10784 8888
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 11238 8848 11244 8900
rect 11296 8848 11302 8900
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 14921 8891 14979 8897
rect 14921 8888 14933 8891
rect 14332 8860 14933 8888
rect 14332 8848 14338 8860
rect 14921 8857 14933 8860
rect 14967 8857 14979 8891
rect 14921 8851 14979 8857
rect 9508 8792 9812 8820
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 11256 8820 11284 8848
rect 10652 8792 11284 8820
rect 10652 8780 10658 8792
rect 12894 8780 12900 8832
rect 12952 8780 12958 8832
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14734 8820 14740 8832
rect 14415 8792 14740 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 1104 8730 16284 8752
rect 1104 8678 3507 8730
rect 3559 8678 3571 8730
rect 3623 8678 3635 8730
rect 3687 8678 3699 8730
rect 3751 8678 3763 8730
rect 3815 8678 7302 8730
rect 7354 8678 7366 8730
rect 7418 8678 7430 8730
rect 7482 8678 7494 8730
rect 7546 8678 7558 8730
rect 7610 8678 11097 8730
rect 11149 8678 11161 8730
rect 11213 8678 11225 8730
rect 11277 8678 11289 8730
rect 11341 8678 11353 8730
rect 11405 8678 14892 8730
rect 14944 8678 14956 8730
rect 15008 8678 15020 8730
rect 15072 8678 15084 8730
rect 15136 8678 15148 8730
rect 15200 8678 16284 8730
rect 1104 8656 16284 8678
rect 6822 8616 6828 8628
rect 6380 8588 6828 8616
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6380 8480 6408 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9306 8616 9312 8628
rect 9263 8588 9312 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10226 8616 10232 8628
rect 10183 8588 10232 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10778 8576 10784 8628
rect 10836 8576 10842 8628
rect 10962 8625 10968 8628
rect 10949 8619 10968 8625
rect 10949 8585 10961 8619
rect 10949 8579 10968 8585
rect 10962 8576 10968 8579
rect 11020 8576 11026 8628
rect 12894 8616 12900 8628
rect 12406 8588 12900 8616
rect 7098 8508 7104 8560
rect 7156 8508 7162 8560
rect 8220 8548 8248 8576
rect 10594 8548 10600 8560
rect 8220 8520 10600 8548
rect 6043 8452 6408 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 9324 8489 9352 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 11149 8551 11207 8557
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 11422 8548 11428 8560
rect 11195 8520 11428 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 8536 8452 8953 8480
rect 8536 8440 8542 8452
rect 8941 8449 8953 8452
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 10192 8452 10333 8480
rect 10192 8440 10198 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5316 8384 6377 8412
rect 5316 8372 5322 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6365 8375 6423 8381
rect 6472 8384 6653 8412
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6472 8344 6500 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10428 8412 10456 8443
rect 10612 8421 10640 8508
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10008 8384 10456 8412
rect 10597 8415 10655 8421
rect 10008 8372 10014 8384
rect 10597 8381 10609 8415
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 6227 8316 6500 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 9214 8344 9220 8356
rect 7800 8316 9220 8344
rect 7800 8304 7806 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 10704 8344 10732 8443
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12406 8480 12434 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13446 8616 13452 8628
rect 13035 8588 13452 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 14274 8576 14280 8628
rect 14332 8576 14338 8628
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 13357 8551 13415 8557
rect 13357 8517 13369 8551
rect 13403 8548 13415 8551
rect 13998 8548 14004 8560
rect 13403 8520 14004 8548
rect 13403 8517 13415 8520
rect 13357 8511 13415 8517
rect 12023 8452 12434 8480
rect 12897 8483 12955 8489
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13372 8480 13400 8511
rect 13998 8508 14004 8520
rect 14056 8508 14062 8560
rect 12943 8452 13400 8480
rect 13909 8483 13967 8489
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14292 8480 14320 8576
rect 13955 8452 14320 8480
rect 14553 8483 14611 8489
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15304 8480 15332 8576
rect 15151 8452 15332 8480
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8412 12403 8415
rect 12802 8412 12808 8424
rect 12391 8384 12808 8412
rect 12391 8381 12403 8384
rect 12345 8375 12403 8381
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 13280 8384 13461 8412
rect 13280 8356 13308 8384
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 14182 8412 14188 8424
rect 13679 8384 14188 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 14182 8372 14188 8384
rect 14240 8412 14246 8424
rect 14277 8415 14335 8421
rect 14277 8412 14289 8415
rect 14240 8384 14289 8412
rect 14240 8372 14246 8384
rect 14277 8381 14289 8384
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8381 14519 8415
rect 14568 8412 14596 8443
rect 15580 8412 15608 8576
rect 14568 8384 15608 8412
rect 14461 8375 14519 8381
rect 13262 8344 13268 8356
rect 10704 8316 13268 8344
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 8386 8236 8392 8288
rect 8444 8236 8450 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 10962 8236 10968 8288
rect 11020 8236 11026 8288
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 12161 8279 12219 8285
rect 12161 8245 12173 8279
rect 12207 8276 12219 8279
rect 12250 8276 12256 8288
rect 12207 8248 12256 8276
rect 12207 8245 12219 8248
rect 12161 8239 12219 8245
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 14090 8236 14096 8288
rect 14148 8236 14154 8288
rect 14292 8276 14320 8375
rect 14476 8344 14504 8375
rect 15838 8344 15844 8356
rect 14476 8316 15844 8344
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 14642 8276 14648 8288
rect 14292 8248 14648 8276
rect 14642 8236 14648 8248
rect 14700 8236 14706 8288
rect 14921 8279 14979 8285
rect 14921 8245 14933 8279
rect 14967 8276 14979 8279
rect 15470 8276 15476 8288
rect 14967 8248 15476 8276
rect 14967 8245 14979 8248
rect 14921 8239 14979 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 1104 8186 16284 8208
rect 1104 8134 2847 8186
rect 2899 8134 2911 8186
rect 2963 8134 2975 8186
rect 3027 8134 3039 8186
rect 3091 8134 3103 8186
rect 3155 8134 6642 8186
rect 6694 8134 6706 8186
rect 6758 8134 6770 8186
rect 6822 8134 6834 8186
rect 6886 8134 6898 8186
rect 6950 8134 10437 8186
rect 10489 8134 10501 8186
rect 10553 8134 10565 8186
rect 10617 8134 10629 8186
rect 10681 8134 10693 8186
rect 10745 8134 14232 8186
rect 14284 8134 14296 8186
rect 14348 8134 14360 8186
rect 14412 8134 14424 8186
rect 14476 8134 14488 8186
rect 14540 8134 16284 8186
rect 1104 8112 16284 8134
rect 8018 8072 8024 8084
rect 4080 8044 8024 8072
rect 2685 8007 2743 8013
rect 2685 7973 2697 8007
rect 2731 7973 2743 8007
rect 2685 7967 2743 7973
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2700 7868 2728 7967
rect 3234 7896 3240 7948
rect 3292 7896 3298 7948
rect 2639 7840 2728 7868
rect 3053 7871 3111 7877
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3970 7868 3976 7880
rect 3099 7840 3976 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3970 7828 3976 7840
rect 4028 7868 4034 7880
rect 4080 7877 4108 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 9180 8044 9229 8072
rect 9180 8032 9186 8044
rect 9217 8041 9229 8044
rect 9263 8072 9275 8075
rect 9490 8072 9496 8084
rect 9263 8044 9496 8072
rect 9263 8041 9275 8044
rect 9217 8035 9275 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10686 8072 10692 8084
rect 9916 8044 10692 8072
rect 9916 8032 9922 8044
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13320 8044 13737 8072
rect 13320 8032 13326 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 14090 8032 14096 8084
rect 14148 8032 14154 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 12250 7896 12256 7948
rect 12308 7896 12314 7948
rect 14108 7936 14136 8032
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 14108 7908 14381 7936
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 4028 7840 4077 7868
rect 4028 7828 4034 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 4065 7831 4123 7837
rect 5276 7840 7113 7868
rect 5276 7812 5304 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 8202 7868 8208 7880
rect 7101 7831 7159 7837
rect 7300 7840 8208 7868
rect 5258 7800 5264 7812
rect 4540 7772 5264 7800
rect 4540 7744 4568 7772
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7300 7800 7328 7840
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 11974 7868 11980 7880
rect 9539 7840 11980 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 7055 7772 7328 7800
rect 7368 7803 7426 7809
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7368 7769 7380 7803
rect 7414 7769 7426 7803
rect 7368 7763 7426 7769
rect 9033 7803 9091 7809
rect 9033 7769 9045 7803
rect 9079 7800 9091 7803
rect 9582 7800 9588 7812
rect 9079 7772 9588 7800
rect 9079 7769 9091 7772
rect 9033 7763 9091 7769
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 3142 7692 3148 7744
rect 3200 7692 3206 7744
rect 4522 7692 4528 7744
rect 4580 7692 4586 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7392 7732 7420 7763
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 9760 7803 9818 7809
rect 9760 7769 9772 7803
rect 9806 7800 9818 7803
rect 11514 7800 11520 7812
rect 9806 7772 11520 7800
rect 9806 7769 9818 7772
rect 9760 7763 9818 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12406 7772 12742 7800
rect 6972 7704 7420 7732
rect 6972 7692 6978 7704
rect 9214 7692 9220 7744
rect 9272 7741 9278 7744
rect 9272 7735 9291 7741
rect 9279 7701 9291 7735
rect 9272 7695 9291 7701
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9858 7732 9864 7744
rect 9447 7704 9864 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9272 7692 9278 7695
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 12406 7732 12434 7772
rect 10744 7704 12434 7732
rect 12636 7732 12664 7772
rect 13814 7732 13820 7744
rect 12636 7704 13820 7732
rect 10744 7692 10750 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 1104 7642 16284 7664
rect 1104 7590 3507 7642
rect 3559 7590 3571 7642
rect 3623 7590 3635 7642
rect 3687 7590 3699 7642
rect 3751 7590 3763 7642
rect 3815 7590 7302 7642
rect 7354 7590 7366 7642
rect 7418 7590 7430 7642
rect 7482 7590 7494 7642
rect 7546 7590 7558 7642
rect 7610 7590 11097 7642
rect 11149 7590 11161 7642
rect 11213 7590 11225 7642
rect 11277 7590 11289 7642
rect 11341 7590 11353 7642
rect 11405 7590 14892 7642
rect 14944 7590 14956 7642
rect 15008 7590 15020 7642
rect 15072 7590 15084 7642
rect 15136 7590 15148 7642
rect 15200 7590 16284 7642
rect 1104 7568 16284 7590
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3200 7500 3893 7528
rect 3200 7488 3206 7500
rect 3881 7497 3893 7500
rect 3927 7497 3939 7531
rect 3881 7491 3939 7497
rect 3970 7488 3976 7540
rect 4028 7488 4034 7540
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7587 7531 7645 7537
rect 7587 7497 7599 7531
rect 7633 7528 7645 7531
rect 7742 7528 7748 7540
rect 7633 7500 7748 7528
rect 7633 7497 7645 7500
rect 7587 7491 7645 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8386 7528 8392 7540
rect 8251 7500 8392 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 2317 7463 2375 7469
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 2424 7460 2452 7488
rect 2363 7432 2452 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 3326 7420 3332 7472
rect 3384 7420 3390 7472
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 1596 7256 1624 7355
rect 1670 7284 1676 7336
rect 1728 7284 1734 7336
rect 2038 7284 2044 7336
rect 2096 7284 2102 7336
rect 3050 7324 3056 7336
rect 2148 7296 3056 7324
rect 2148 7256 2176 7296
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 3988 7324 4016 7488
rect 5994 7420 6000 7472
rect 6052 7460 6058 7472
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 6052 7432 7389 7460
rect 6052 7420 6058 7432
rect 7377 7429 7389 7432
rect 7423 7429 7435 7463
rect 7377 7423 7435 7429
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7852 7392 7880 7491
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9398 7528 9404 7540
rect 9171 7500 9404 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 9950 7528 9956 7540
rect 9631 7500 9956 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 12802 7488 12808 7540
rect 12860 7488 12866 7540
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 12952 7500 13952 7528
rect 12952 7488 12958 7500
rect 10720 7463 10778 7469
rect 10720 7429 10732 7463
rect 10766 7460 10778 7463
rect 11238 7460 11244 7472
rect 10766 7432 11244 7460
rect 10766 7429 10778 7432
rect 10720 7423 10778 7429
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 13924 7460 13952 7500
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14056 7500 14688 7528
rect 14056 7488 14062 7500
rect 14660 7460 14688 7500
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14792 7500 15025 7528
rect 14792 7488 14798 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 15105 7463 15163 7469
rect 15105 7460 15117 7463
rect 13846 7432 14596 7460
rect 14660 7432 15117 7460
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 6779 7364 7880 7392
rect 8312 7364 9045 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 3835 7296 4016 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4430 7284 4436 7336
rect 4488 7324 4494 7336
rect 4632 7324 4660 7355
rect 4488 7296 4660 7324
rect 4488 7284 4494 7296
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 8312 7333 8340 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11974 7392 11980 7404
rect 11011 7364 11980 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 14568 7392 14596 7432
rect 15105 7429 15117 7432
rect 15151 7429 15163 7463
rect 15105 7423 15163 7429
rect 15396 7392 15424 7488
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 14568 7364 15332 7392
rect 15396 7364 15669 7392
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 7248 7296 8309 7324
rect 7248 7284 7254 7296
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 1596 7228 2176 7256
rect 7745 7259 7803 7265
rect 7745 7225 7757 7259
rect 7791 7256 7803 7259
rect 8404 7256 8432 7287
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13964 7296 14289 7324
rect 13964 7284 13970 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7293 14611 7327
rect 14553 7287 14611 7293
rect 7791 7228 8432 7256
rect 9493 7259 9551 7265
rect 7791 7225 7803 7228
rect 7745 7219 7803 7225
rect 9493 7225 9505 7259
rect 9539 7256 9551 7259
rect 9539 7228 10088 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 1946 7148 1952 7200
rect 2004 7148 2010 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7561 7191 7619 7197
rect 7561 7188 7573 7191
rect 7064 7160 7573 7188
rect 7064 7148 7070 7160
rect 7561 7157 7573 7160
rect 7607 7188 7619 7191
rect 9398 7188 9404 7200
rect 7607 7160 9404 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 10060 7188 10088 7228
rect 11146 7188 11152 7200
rect 10060 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14568 7188 14596 7287
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14700 7296 15209 7324
rect 14700 7284 14706 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15304 7324 15332 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15378 7324 15384 7336
rect 15304 7296 15384 7324
rect 15197 7287 15255 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 14148 7160 14596 7188
rect 14148 7148 14154 7160
rect 14642 7148 14648 7200
rect 14700 7148 14706 7200
rect 15470 7148 15476 7200
rect 15528 7148 15534 7200
rect 1104 7098 16284 7120
rect 1104 7046 2847 7098
rect 2899 7046 2911 7098
rect 2963 7046 2975 7098
rect 3027 7046 3039 7098
rect 3091 7046 3103 7098
rect 3155 7046 6642 7098
rect 6694 7046 6706 7098
rect 6758 7046 6770 7098
rect 6822 7046 6834 7098
rect 6886 7046 6898 7098
rect 6950 7046 10437 7098
rect 10489 7046 10501 7098
rect 10553 7046 10565 7098
rect 10617 7046 10629 7098
rect 10681 7046 10693 7098
rect 10745 7046 14232 7098
rect 14284 7046 14296 7098
rect 14348 7046 14360 7098
rect 14412 7046 14424 7098
rect 14476 7046 14488 7098
rect 14540 7046 16284 7098
rect 1104 7024 16284 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2114 6987 2172 6993
rect 2114 6984 2126 6987
rect 2004 6956 2126 6984
rect 2004 6944 2010 6956
rect 2114 6953 2126 6956
rect 2160 6953 2172 6987
rect 2114 6947 2172 6953
rect 11238 6944 11244 6996
rect 11296 6944 11302 6996
rect 13541 6987 13599 6993
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 13906 6984 13912 6996
rect 13587 6956 13912 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 14356 6987 14414 6993
rect 14356 6953 14368 6987
rect 14402 6984 14414 6987
rect 15470 6984 15476 6996
rect 14402 6956 15476 6984
rect 14402 6953 14414 6956
rect 14356 6947 14414 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 3326 6808 3332 6860
rect 3384 6808 3390 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6848 6423 6851
rect 6546 6848 6552 6860
rect 6411 6820 6552 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6848 9827 6851
rect 9858 6848 9864 6860
rect 9815 6820 9864 6848
rect 9815 6817 9827 6820
rect 9769 6811 9827 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10928 6820 11069 6848
rect 10928 6808 10934 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 14090 6848 14096 6860
rect 12032 6820 14096 6848
rect 12032 6808 12038 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 3344 6780 3372 6808
rect 3266 6752 3372 6780
rect 1857 6743 1915 6749
rect 1872 6712 1900 6743
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 1872 6684 2084 6712
rect 2056 6656 2084 6684
rect 6472 6656 6500 6743
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11204 6752 11437 6780
rect 11204 6740 11210 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 7190 6672 7196 6724
rect 7248 6672 7254 6724
rect 9953 6715 10011 6721
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 10505 6715 10563 6721
rect 10505 6712 10517 6715
rect 9999 6684 10517 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 10505 6681 10517 6684
rect 10551 6681 10563 6715
rect 10505 6675 10563 6681
rect 2038 6604 2044 6656
rect 2096 6604 2102 6656
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3476 6616 3617 6644
rect 3476 6604 3482 6616
rect 3605 6613 3617 6616
rect 3651 6644 3663 6647
rect 4430 6644 4436 6656
rect 3651 6616 4436 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 6454 6604 6460 6656
rect 6512 6604 6518 6656
rect 7208 6644 7236 6672
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 7208 6616 9873 6644
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 9861 6607 9919 6613
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6644 10379 6647
rect 11698 6644 11704 6656
rect 10367 6616 11704 6644
rect 10367 6613 10379 6616
rect 10321 6607 10379 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 13372 6644 13400 6743
rect 15378 6740 15384 6792
rect 15436 6780 15442 6792
rect 15436 6752 15502 6780
rect 15436 6740 15442 6752
rect 14642 6672 14648 6724
rect 14700 6672 14706 6724
rect 14660 6644 14688 6672
rect 13372 6616 14688 6644
rect 15838 6604 15844 6656
rect 15896 6604 15902 6656
rect 1104 6554 16284 6576
rect 1104 6502 3507 6554
rect 3559 6502 3571 6554
rect 3623 6502 3635 6554
rect 3687 6502 3699 6554
rect 3751 6502 3763 6554
rect 3815 6502 7302 6554
rect 7354 6502 7366 6554
rect 7418 6502 7430 6554
rect 7482 6502 7494 6554
rect 7546 6502 7558 6554
rect 7610 6502 11097 6554
rect 11149 6502 11161 6554
rect 11213 6502 11225 6554
rect 11277 6502 11289 6554
rect 11341 6502 11353 6554
rect 11405 6502 14892 6554
rect 14944 6502 14956 6554
rect 15008 6502 15020 6554
rect 15072 6502 15084 6554
rect 15136 6502 15148 6554
rect 15200 6502 16284 6554
rect 1104 6480 16284 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 1728 6412 2697 6440
rect 1728 6400 1734 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 3326 6400 3332 6452
rect 3384 6400 3390 6452
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8996 6412 9505 6440
rect 8996 6400 9002 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10962 6440 10968 6452
rect 9907 6412 10968 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15654 6440 15660 6452
rect 15243 6412 15660 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 3344 6372 3372 6400
rect 3344 6344 5198 6372
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 9272 6344 9689 6372
rect 9272 6332 9278 6344
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 9677 6335 9735 6341
rect 10045 6375 10103 6381
rect 10045 6341 10057 6375
rect 10091 6372 10103 6375
rect 10134 6372 10140 6384
rect 10091 6344 10140 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10134 6332 10140 6344
rect 10192 6372 10198 6384
rect 11422 6372 11428 6384
rect 10192 6344 11428 6372
rect 10192 6332 10198 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 3418 6304 3424 6316
rect 3375 6276 3424 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6932 6276 7113 6304
rect 2056 6236 2084 6264
rect 4430 6236 4436 6248
rect 2056 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4706 6196 4712 6248
rect 4764 6196 4770 6248
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6454 6236 6460 6248
rect 6227 6208 6460 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6454 6196 6460 6208
rect 6512 6236 6518 6248
rect 6932 6245 6960 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 7101 6267 7159 6273
rect 9692 6276 9781 6304
rect 9692 6248 9720 6276
rect 9769 6273 9781 6276
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10008 6276 10793 6304
rect 10008 6264 10014 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6512 6208 6929 6236
rect 6512 6196 6518 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 9674 6196 9680 6248
rect 9732 6196 9738 6248
rect 9766 6128 9772 6180
rect 9824 6128 9830 6180
rect 6362 6060 6368 6112
rect 6420 6060 6426 6112
rect 9784 6100 9812 6128
rect 10870 6100 10876 6112
rect 9784 6072 10876 6100
rect 10870 6060 10876 6072
rect 10928 6100 10934 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10928 6072 10977 6100
rect 10928 6060 10934 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 1104 6010 16284 6032
rect 1104 5958 2847 6010
rect 2899 5958 2911 6010
rect 2963 5958 2975 6010
rect 3027 5958 3039 6010
rect 3091 5958 3103 6010
rect 3155 5958 6642 6010
rect 6694 5958 6706 6010
rect 6758 5958 6770 6010
rect 6822 5958 6834 6010
rect 6886 5958 6898 6010
rect 6950 5958 10437 6010
rect 10489 5958 10501 6010
rect 10553 5958 10565 6010
rect 10617 5958 10629 6010
rect 10681 5958 10693 6010
rect 10745 5958 14232 6010
rect 14284 5958 14296 6010
rect 14348 5958 14360 6010
rect 14412 5958 14424 6010
rect 14476 5958 14488 6010
rect 14540 5958 16284 6010
rect 1104 5936 16284 5958
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 4764 5868 5181 5896
rect 4764 5856 4770 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 5169 5859 5227 5865
rect 6362 5856 6368 5908
rect 6420 5856 6426 5908
rect 10134 5896 10140 5908
rect 9692 5868 10140 5896
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5810 5760 5816 5772
rect 5675 5732 5816 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5810 5720 5816 5732
rect 5868 5760 5874 5772
rect 6270 5760 6276 5772
rect 5868 5732 6276 5760
rect 5868 5720 5874 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 6380 5692 6408 5856
rect 7190 5788 7196 5840
rect 7248 5788 7254 5840
rect 6730 5720 6736 5772
rect 6788 5720 6794 5772
rect 9692 5760 9720 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 11974 5896 11980 5908
rect 11931 5868 11980 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15289 5899 15347 5905
rect 15289 5896 15301 5899
rect 14792 5868 15301 5896
rect 14792 5856 14798 5868
rect 15289 5865 15301 5868
rect 15335 5865 15347 5899
rect 15289 5859 15347 5865
rect 15838 5856 15844 5908
rect 15896 5856 15902 5908
rect 15856 5769 15884 5856
rect 15841 5763 15899 5769
rect 9684 5732 9720 5760
rect 10244 5732 11008 5760
rect 9684 5711 9712 5732
rect 9653 5705 9712 5711
rect 5583 5664 6408 5692
rect 6825 5695 6883 5701
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 7190 5692 7196 5704
rect 6871 5664 7196 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9653 5671 9665 5705
rect 9699 5674 9712 5705
rect 9699 5671 9711 5674
rect 9653 5665 9711 5671
rect 9757 5652 9763 5704
rect 9815 5652 9821 5704
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 9508 5624 9536 5652
rect 9759 5639 9771 5652
rect 9805 5639 9817 5652
rect 9759 5633 9817 5639
rect 9508 5596 9720 5624
rect 9582 5516 9588 5568
rect 9640 5516 9646 5568
rect 9692 5556 9720 5596
rect 9876 5556 9904 5655
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10145 5695 10203 5701
rect 10145 5661 10157 5695
rect 10191 5692 10203 5695
rect 10244 5692 10272 5732
rect 10980 5704 11008 5732
rect 15841 5729 15853 5763
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 10191 5664 10272 5692
rect 10191 5661 10203 5664
rect 10145 5655 10203 5661
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10376 5664 10425 5692
rect 10376 5652 10382 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 9692 5528 9904 5556
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 12066 5556 12072 5568
rect 10367 5528 12072 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 1104 5466 16284 5488
rect 1104 5414 3507 5466
rect 3559 5414 3571 5466
rect 3623 5414 3635 5466
rect 3687 5414 3699 5466
rect 3751 5414 3763 5466
rect 3815 5414 7302 5466
rect 7354 5414 7366 5466
rect 7418 5414 7430 5466
rect 7482 5414 7494 5466
rect 7546 5414 7558 5466
rect 7610 5414 11097 5466
rect 11149 5414 11161 5466
rect 11213 5414 11225 5466
rect 11277 5414 11289 5466
rect 11341 5414 11353 5466
rect 11405 5414 14892 5466
rect 14944 5414 14956 5466
rect 15008 5414 15020 5466
rect 15072 5414 15084 5466
rect 15136 5414 15148 5466
rect 15200 5414 16284 5466
rect 1104 5392 16284 5414
rect 5810 5352 5816 5364
rect 5552 5324 5816 5352
rect 2869 5287 2927 5293
rect 2869 5253 2881 5287
rect 2915 5284 2927 5287
rect 3234 5284 3240 5296
rect 2915 5256 3240 5284
rect 2915 5253 2927 5256
rect 2869 5247 2927 5253
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 5552 5225 5580 5324
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9582 5352 9588 5364
rect 9088 5324 9588 5352
rect 9088 5312 9094 5324
rect 9582 5312 9588 5324
rect 9640 5352 9646 5364
rect 10042 5352 10048 5364
rect 9640 5324 10048 5352
rect 9640 5312 9646 5324
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 6457 5287 6515 5293
rect 6457 5284 6469 5287
rect 5736 5256 6469 5284
rect 5736 5225 5764 5256
rect 6457 5253 6469 5256
rect 6503 5253 6515 5287
rect 9950 5284 9956 5296
rect 6457 5247 6515 5253
rect 7484 5256 9956 5284
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2280 5188 2697 5216
rect 2280 5176 2286 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5868 5188 6009 5216
rect 5868 5176 5874 5188
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6043 5188 6377 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6595 5188 6837 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6730 5148 6736 5160
rect 6227 5120 6736 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6730 5108 6736 5120
rect 6788 5148 6794 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6788 5120 7389 5148
rect 6788 5108 6794 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 7484 5080 7512 5256
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9582 5216 9588 5228
rect 9456 5188 9588 5216
rect 9456 5176 9462 5188
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 10060 5157 10088 5312
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11388 5256 12296 5284
rect 11388 5244 11394 5256
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 12268 5225 12296 5256
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10091 5120 10272 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 9968 5080 9996 5111
rect 10134 5080 10140 5092
rect 5224 5052 7512 5080
rect 8680 5052 9904 5080
rect 9968 5052 10140 5080
rect 5224 5040 5230 5052
rect 8680 5024 8708 5052
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 4154 5012 4160 5024
rect 3099 4984 4160 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5684 4984 5733 5012
rect 5684 4972 5690 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 9876 5012 9904 5052
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 10244 5080 10272 5120
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5148 10839 5151
rect 10962 5148 10968 5160
rect 10827 5120 10968 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12360 5148 12388 5179
rect 11388 5120 12388 5148
rect 11388 5108 11394 5120
rect 12544 5080 12572 5179
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 10244 5052 12572 5080
rect 10410 5012 10416 5024
rect 9876 4984 10416 5012
rect 9769 4975 9827 4981
rect 10410 4972 10416 4984
rect 10468 5012 10474 5024
rect 10778 5012 10784 5024
rect 10468 4984 10784 5012
rect 10468 4972 10474 4984
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 12802 4972 12808 5024
rect 12860 4972 12866 5024
rect 1104 4922 16284 4944
rect 1104 4870 2847 4922
rect 2899 4870 2911 4922
rect 2963 4870 2975 4922
rect 3027 4870 3039 4922
rect 3091 4870 3103 4922
rect 3155 4870 6642 4922
rect 6694 4870 6706 4922
rect 6758 4870 6770 4922
rect 6822 4870 6834 4922
rect 6886 4870 6898 4922
rect 6950 4870 10437 4922
rect 10489 4870 10501 4922
rect 10553 4870 10565 4922
rect 10617 4870 10629 4922
rect 10681 4870 10693 4922
rect 10745 4870 14232 4922
rect 14284 4870 14296 4922
rect 14348 4870 14360 4922
rect 14412 4870 14424 4922
rect 14476 4870 14488 4922
rect 14540 4870 16284 4922
rect 1104 4848 16284 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3326 4808 3332 4820
rect 3283 4780 3332 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 4430 4768 4436 4820
rect 4488 4768 4494 4820
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6604 4780 7021 4808
rect 6604 4768 6610 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 2682 4700 2688 4752
rect 2740 4700 2746 4752
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 2700 4672 2728 4700
rect 2639 4644 2728 4672
rect 3344 4672 3372 4768
rect 4448 4740 4476 4768
rect 4448 4712 5304 4740
rect 5276 4684 5304 4712
rect 3344 4644 4476 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 2731 4576 3801 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 2240 4536 2268 4567
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4304 4576 4353 4604
rect 4304 4564 4310 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 3234 4536 3240 4548
rect 2240 4508 3240 4536
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 3329 4539 3387 4545
rect 3329 4505 3341 4539
rect 3375 4505 3387 4539
rect 4448 4536 4476 4644
rect 5258 4632 5264 4684
rect 5316 4632 5322 4684
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5626 4672 5632 4684
rect 5583 4644 5632 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 5166 4604 5172 4616
rect 4580 4576 5172 4604
rect 4580 4564 4586 4576
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 7024 4604 7052 4771
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7248 4780 7297 4808
rect 7248 4768 7254 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 8662 4768 8668 4820
rect 8720 4768 8726 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 9048 4780 10885 4808
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7024 4576 7573 4604
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 9048 4604 9076 4780
rect 10873 4777 10885 4780
rect 10919 4808 10931 4811
rect 10962 4808 10968 4820
rect 10919 4780 10968 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11228 4811 11286 4817
rect 11228 4777 11240 4811
rect 11274 4808 11286 4811
rect 11422 4808 11428 4820
rect 11274 4780 11428 4808
rect 11274 4777 11286 4780
rect 11228 4771 11286 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 9180 4644 10977 4672
rect 9180 4632 9186 4644
rect 10965 4641 10977 4644
rect 11011 4672 11023 4675
rect 11974 4672 11980 4684
rect 11011 4644 11980 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12894 4604 12900 4616
rect 8803 4576 9076 4604
rect 12406 4576 12900 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 5994 4536 6000 4548
rect 4448 4508 5212 4536
rect 3329 4499 3387 4505
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 2004 4440 2053 4468
rect 2004 4428 2010 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 2041 4431 2099 4437
rect 2314 4428 2320 4480
rect 2372 4428 2378 4480
rect 3344 4468 3372 4499
rect 4338 4468 4344 4480
rect 3344 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4468 4402 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 4396 4440 4721 4468
rect 4396 4428 4402 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 5184 4468 5212 4508
rect 5552 4508 6000 4536
rect 5552 4468 5580 4508
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 7469 4539 7527 4545
rect 7469 4505 7481 4539
rect 7515 4536 7527 4539
rect 8202 4536 8208 4548
rect 7515 4508 8208 4536
rect 7515 4505 7527 4508
rect 7469 4499 7527 4505
rect 8202 4496 8208 4508
rect 8260 4536 8266 4548
rect 8588 4536 8616 4567
rect 8260 4508 8616 4536
rect 9401 4539 9459 4545
rect 8260 4496 8266 4508
rect 9401 4505 9413 4539
rect 9447 4505 9459 4539
rect 9401 4499 9459 4505
rect 5184 4440 5580 4468
rect 4709 4431 4767 4437
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 5776 4440 7113 4468
rect 5776 4428 5782 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 7269 4471 7327 4477
rect 7269 4437 7281 4471
rect 7315 4468 7327 4471
rect 8110 4468 8116 4480
rect 7315 4440 8116 4468
rect 7315 4437 7327 4440
rect 7269 4431 7327 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 9416 4468 9444 4499
rect 9858 4496 9864 4548
rect 9916 4496 9922 4548
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 10836 4508 11730 4536
rect 10836 4496 10842 4508
rect 9272 4440 9444 4468
rect 9272 4428 9278 4440
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 11330 4468 11336 4480
rect 9640 4440 11336 4468
rect 9640 4428 9646 4440
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 11624 4468 11652 4508
rect 12406 4468 12434 4576
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 11624 4440 12434 4468
rect 12710 4428 12716 4480
rect 12768 4428 12774 4480
rect 1104 4378 16284 4400
rect 1104 4326 3507 4378
rect 3559 4326 3571 4378
rect 3623 4326 3635 4378
rect 3687 4326 3699 4378
rect 3751 4326 3763 4378
rect 3815 4326 7302 4378
rect 7354 4326 7366 4378
rect 7418 4326 7430 4378
rect 7482 4326 7494 4378
rect 7546 4326 7558 4378
rect 7610 4326 11097 4378
rect 11149 4326 11161 4378
rect 11213 4326 11225 4378
rect 11277 4326 11289 4378
rect 11341 4326 11353 4378
rect 11405 4326 14892 4378
rect 14944 4326 14956 4378
rect 15008 4326 15020 4378
rect 15072 4326 15084 4378
rect 15136 4326 15148 4378
rect 15200 4326 16284 4378
rect 1104 4304 16284 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3292 4236 3893 4264
rect 3292 4224 3298 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 3881 4227 3939 4233
rect 9030 4224 9036 4276
rect 9088 4224 9094 4276
rect 9122 4224 9128 4276
rect 9180 4224 9186 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 10778 4264 10784 4276
rect 9916 4236 10784 4264
rect 9916 4224 9922 4236
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 2222 4196 2228 4208
rect 1964 4168 2228 4196
rect 1964 4137 1992 4168
rect 2222 4156 2228 4168
rect 2280 4156 2286 4208
rect 2314 4156 2320 4208
rect 2372 4156 2378 4208
rect 3326 4156 3332 4208
rect 3384 4156 3390 4208
rect 6181 4199 6239 4205
rect 5828 4168 6132 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 1780 3924 1808 4091
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2682 4060 2688 4072
rect 1903 4032 2688 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2682 4020 2688 4032
rect 2740 4060 2746 4072
rect 4080 4060 4108 4091
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 5718 4128 5724 4140
rect 5675 4100 5724 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 5828 4137 5856 4168
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5902 4088 5908 4140
rect 5960 4088 5966 4140
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6104 4128 6132 4168
rect 6181 4165 6193 4199
rect 6227 4196 6239 4199
rect 7561 4199 7619 4205
rect 7561 4196 7573 4199
rect 6227 4168 7573 4196
rect 6227 4165 6239 4168
rect 6181 4159 6239 4165
rect 7561 4165 7573 4168
rect 7607 4165 7619 4199
rect 9140 4196 9168 4224
rect 9876 4196 9904 4224
rect 9140 4168 9260 4196
rect 9876 4168 9982 4196
rect 7561 4159 7619 4165
rect 6104 4100 6224 4128
rect 5997 4091 6055 4097
rect 2740 4032 4108 4060
rect 2740 4020 2746 4032
rect 4246 4020 4252 4072
rect 4304 4020 4310 4072
rect 6012 4060 6040 4091
rect 6086 4060 6092 4072
rect 5736 4032 6092 4060
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 4264 3992 4292 4020
rect 3835 3964 4292 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 3050 3924 3056 3936
rect 1780 3896 3056 3924
rect 3050 3884 3056 3896
rect 3108 3924 3114 3936
rect 3970 3924 3976 3936
rect 3108 3896 3976 3924
rect 3108 3884 3114 3896
rect 3970 3884 3976 3896
rect 4028 3924 4034 3936
rect 5736 3924 5764 4032
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6196 4001 6224 4100
rect 7190 4088 7196 4140
rect 7248 4088 7254 4140
rect 8110 4088 8116 4140
rect 8168 4088 8174 4140
rect 9232 4137 9260 4168
rect 12894 4156 12900 4208
rect 12952 4156 12958 4208
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 9674 4128 9680 4140
rect 9631 4100 9680 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 7208 4060 7236 4088
rect 8312 4060 8340 4091
rect 7208 4032 8340 4060
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 4028 3896 5764 3924
rect 4028 3884 4034 3896
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5960 3896 6561 3924
rect 5960 3884 5966 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 8662 3884 8668 3936
rect 8720 3884 8726 3936
rect 8864 3924 8892 4091
rect 9140 4060 9168 4091
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 11974 4128 11980 4140
rect 11563 4100 11980 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 13311 4131 13369 4137
rect 13311 4097 13323 4131
rect 13357 4128 13369 4131
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13357 4100 13461 4128
rect 13357 4097 13369 4100
rect 13311 4091 13369 4097
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 9490 4060 9496 4072
rect 9140 4032 9496 4060
rect 9490 4020 9496 4032
rect 9548 4060 9554 4072
rect 11054 4060 11060 4072
rect 9548 4032 11060 4060
rect 9548 4020 9554 4032
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 12802 4060 12808 4072
rect 11931 4032 12808 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 11422 3992 11428 4004
rect 10336 3964 11428 3992
rect 9766 3924 9772 3936
rect 8864 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3924 9830 3936
rect 10336 3924 10364 3964
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 9824 3896 10364 3924
rect 11011 3927 11069 3933
rect 9824 3884 9830 3896
rect 11011 3893 11023 3927
rect 11057 3924 11069 3927
rect 12618 3924 12624 3936
rect 11057 3896 12624 3924
rect 11057 3893 11069 3896
rect 11011 3887 11069 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 1104 3834 16284 3856
rect 1104 3782 2847 3834
rect 2899 3782 2911 3834
rect 2963 3782 2975 3834
rect 3027 3782 3039 3834
rect 3091 3782 3103 3834
rect 3155 3782 6642 3834
rect 6694 3782 6706 3834
rect 6758 3782 6770 3834
rect 6822 3782 6834 3834
rect 6886 3782 6898 3834
rect 6950 3782 10437 3834
rect 10489 3782 10501 3834
rect 10553 3782 10565 3834
rect 10617 3782 10629 3834
rect 10681 3782 10693 3834
rect 10745 3782 14232 3834
rect 14284 3782 14296 3834
rect 14348 3782 14360 3834
rect 14412 3782 14424 3834
rect 14476 3782 14488 3834
rect 14540 3782 16284 3834
rect 1104 3760 16284 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 2280 3692 3525 3720
rect 2280 3680 2286 3692
rect 3513 3689 3525 3692
rect 3559 3720 3571 3723
rect 4338 3720 4344 3732
rect 3559 3692 4344 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 5902 3720 5908 3732
rect 5460 3692 5908 3720
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2038 3584 2044 3596
rect 1811 3556 2044 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 5460 3593 5488 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 6144 3692 7144 3720
rect 6144 3680 6150 3692
rect 7116 3652 7144 3692
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7248 3692 7573 3720
rect 7248 3680 7254 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 8662 3680 8668 3732
rect 8720 3680 8726 3732
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10192 3692 11008 3720
rect 10192 3680 10198 3692
rect 8389 3655 8447 3661
rect 8389 3652 8401 3655
rect 7116 3624 8401 3652
rect 8389 3621 8401 3624
rect 8435 3621 8447 3655
rect 8680 3652 8708 3680
rect 10980 3652 11008 3692
rect 11054 3680 11060 3732
rect 11112 3680 11118 3732
rect 12618 3680 12624 3732
rect 12676 3680 12682 3732
rect 11793 3655 11851 3661
rect 11793 3652 11805 3655
rect 8680 3624 9352 3652
rect 10980 3624 11805 3652
rect 8389 3615 8447 3621
rect 5445 3587 5503 3593
rect 3988 3556 5396 3584
rect 3988 3528 4016 3556
rect 3326 3516 3332 3528
rect 3174 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4246 3516 4252 3528
rect 4111 3488 4252 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 5258 3476 5264 3528
rect 5316 3476 5322 3528
rect 5368 3525 5396 3556
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5767 3556 6101 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8110 3516 8116 3528
rect 8067 3488 8116 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2041 3451 2099 3457
rect 2041 3448 2053 3451
rect 2004 3420 2053 3448
rect 2004 3408 2010 3420
rect 2041 3417 2053 3420
rect 2087 3417 2099 3451
rect 5276 3448 5304 3476
rect 5718 3448 5724 3460
rect 5276 3420 5724 3448
rect 2041 3411 2099 3417
rect 5718 3408 5724 3420
rect 5776 3448 5782 3460
rect 5828 3448 5856 3479
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8202 3476 8208 3528
rect 8260 3476 8266 3528
rect 5776 3420 5856 3448
rect 5776 3408 5782 3420
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 8404 3448 8432 3615
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 9180 3556 9229 3584
rect 9180 3544 9186 3556
rect 9217 3553 9229 3556
rect 9263 3553 9275 3587
rect 9324 3584 9352 3624
rect 11793 3621 11805 3624
rect 11839 3621 11851 3655
rect 11793 3615 11851 3621
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9324 3556 9505 3584
rect 9217 3547 9275 3553
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10042 3584 10048 3596
rect 9640 3556 10048 3584
rect 9640 3544 9646 3556
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 11020 3556 11621 3584
rect 11020 3544 11026 3556
rect 11609 3553 11621 3556
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12636 3584 12664 3680
rect 12483 3556 12664 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12710 3516 12716 3528
rect 12667 3488 12716 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 9582 3448 9588 3460
rect 6052 3420 6578 3448
rect 8404 3420 9588 3448
rect 6052 3408 6058 3420
rect 6472 3380 6500 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 9876 3420 9982 3448
rect 9876 3392 9904 3420
rect 6730 3380 6736 3392
rect 6472 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 9858 3340 9864 3392
rect 9916 3340 9922 3392
rect 1104 3290 16284 3312
rect 1104 3238 3507 3290
rect 3559 3238 3571 3290
rect 3623 3238 3635 3290
rect 3687 3238 3699 3290
rect 3751 3238 3763 3290
rect 3815 3238 7302 3290
rect 7354 3238 7366 3290
rect 7418 3238 7430 3290
rect 7482 3238 7494 3290
rect 7546 3238 7558 3290
rect 7610 3238 11097 3290
rect 11149 3238 11161 3290
rect 11213 3238 11225 3290
rect 11277 3238 11289 3290
rect 11341 3238 11353 3290
rect 11405 3238 14892 3290
rect 14944 3238 14956 3290
rect 15008 3238 15020 3290
rect 15072 3238 15084 3290
rect 15136 3238 15148 3290
rect 15200 3238 16284 3290
rect 1104 3216 16284 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5868 3148 6684 3176
rect 5868 3136 5874 3148
rect 6656 3117 6684 3148
rect 8110 3136 8116 3188
rect 8168 3136 8174 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 9916 3148 10701 3176
rect 9916 3136 9922 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 10962 3136 10968 3188
rect 11020 3136 11026 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11480 3148 11621 3176
rect 11480 3136 11486 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 6641 3111 6699 3117
rect 6641 3077 6653 3111
rect 6687 3077 6699 3111
rect 6641 3071 6699 3077
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 9692 3108 9720 3136
rect 10137 3111 10195 3117
rect 10137 3108 10149 3111
rect 6788 3080 7130 3108
rect 9692 3080 10149 3108
rect 6788 3068 6794 3080
rect 10137 3077 10149 3080
rect 10183 3077 10195 3111
rect 10980 3108 11008 3136
rect 10137 3071 10195 3077
rect 10336 3080 11008 3108
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5776 3012 6377 3040
rect 5776 3000 5782 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 8202 3000 8208 3052
rect 8260 3000 8266 3052
rect 10336 3049 10364 3080
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10928 3012 10977 3040
rect 10928 3000 10934 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 12618 3040 12624 3052
rect 11839 3012 12624 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 8220 2972 8248 3000
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 8220 2944 10517 2972
rect 10505 2941 10517 2944
rect 10551 2972 10563 2975
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 10551 2944 11989 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 11977 2941 11989 2944
rect 12023 2972 12035 2975
rect 13814 2972 13820 2984
rect 12023 2944 13820 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 1104 2746 16284 2768
rect 1104 2694 2847 2746
rect 2899 2694 2911 2746
rect 2963 2694 2975 2746
rect 3027 2694 3039 2746
rect 3091 2694 3103 2746
rect 3155 2694 6642 2746
rect 6694 2694 6706 2746
rect 6758 2694 6770 2746
rect 6822 2694 6834 2746
rect 6886 2694 6898 2746
rect 6950 2694 10437 2746
rect 10489 2694 10501 2746
rect 10553 2694 10565 2746
rect 10617 2694 10629 2746
rect 10681 2694 10693 2746
rect 10745 2694 14232 2746
rect 14284 2694 14296 2746
rect 14348 2694 14360 2746
rect 14412 2694 14424 2746
rect 14476 2694 14488 2746
rect 14540 2694 16284 2746
rect 1104 2672 16284 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 4430 2632 4436 2644
rect 1627 2604 4436 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14369 2499 14427 2505
rect 14369 2496 14381 2499
rect 13872 2468 14381 2496
rect 13872 2456 13878 2468
rect 14369 2465 14381 2468
rect 14415 2465 14427 2499
rect 14369 2459 14427 2465
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 1104 2202 16284 2224
rect 1104 2150 3507 2202
rect 3559 2150 3571 2202
rect 3623 2150 3635 2202
rect 3687 2150 3699 2202
rect 3751 2150 3763 2202
rect 3815 2150 7302 2202
rect 7354 2150 7366 2202
rect 7418 2150 7430 2202
rect 7482 2150 7494 2202
rect 7546 2150 7558 2202
rect 7610 2150 11097 2202
rect 11149 2150 11161 2202
rect 11213 2150 11225 2202
rect 11277 2150 11289 2202
rect 11341 2150 11353 2202
rect 11405 2150 14892 2202
rect 14944 2150 14956 2202
rect 15008 2150 15020 2202
rect 15072 2150 15084 2202
rect 15136 2150 15148 2202
rect 15200 2150 16284 2202
rect 1104 2128 16284 2150
<< via1 >>
rect 2847 16838 2899 16890
rect 2911 16838 2963 16890
rect 2975 16838 3027 16890
rect 3039 16838 3091 16890
rect 3103 16838 3155 16890
rect 6642 16838 6694 16890
rect 6706 16838 6758 16890
rect 6770 16838 6822 16890
rect 6834 16838 6886 16890
rect 6898 16838 6950 16890
rect 10437 16838 10489 16890
rect 10501 16838 10553 16890
rect 10565 16838 10617 16890
rect 10629 16838 10681 16890
rect 10693 16838 10745 16890
rect 14232 16838 14284 16890
rect 14296 16838 14348 16890
rect 14360 16838 14412 16890
rect 14424 16838 14476 16890
rect 14488 16838 14540 16890
rect 10232 16600 10284 16652
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 3507 16294 3559 16346
rect 3571 16294 3623 16346
rect 3635 16294 3687 16346
rect 3699 16294 3751 16346
rect 3763 16294 3815 16346
rect 7302 16294 7354 16346
rect 7366 16294 7418 16346
rect 7430 16294 7482 16346
rect 7494 16294 7546 16346
rect 7558 16294 7610 16346
rect 11097 16294 11149 16346
rect 11161 16294 11213 16346
rect 11225 16294 11277 16346
rect 11289 16294 11341 16346
rect 11353 16294 11405 16346
rect 14892 16294 14944 16346
rect 14956 16294 15008 16346
rect 15020 16294 15072 16346
rect 15084 16294 15136 16346
rect 15148 16294 15200 16346
rect 6460 16056 6512 16108
rect 4344 15988 4396 16040
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 6368 15988 6420 16040
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 11612 15988 11664 16040
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 4804 15852 4856 15904
rect 6184 15852 6236 15904
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 9864 15852 9916 15904
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 2847 15750 2899 15802
rect 2911 15750 2963 15802
rect 2975 15750 3027 15802
rect 3039 15750 3091 15802
rect 3103 15750 3155 15802
rect 6642 15750 6694 15802
rect 6706 15750 6758 15802
rect 6770 15750 6822 15802
rect 6834 15750 6886 15802
rect 6898 15750 6950 15802
rect 10437 15750 10489 15802
rect 10501 15750 10553 15802
rect 10565 15750 10617 15802
rect 10629 15750 10681 15802
rect 10693 15750 10745 15802
rect 14232 15750 14284 15802
rect 14296 15750 14348 15802
rect 14360 15750 14412 15802
rect 14424 15750 14476 15802
rect 14488 15750 14540 15802
rect 6184 15648 6236 15700
rect 7380 15648 7432 15700
rect 9036 15648 9088 15700
rect 9588 15648 9640 15700
rect 4528 15512 4580 15564
rect 6184 15512 6236 15564
rect 11520 15580 11572 15632
rect 11796 15580 11848 15632
rect 3976 15444 4028 15496
rect 4252 15444 4304 15496
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 8484 15444 8536 15496
rect 1768 15419 1820 15428
rect 1768 15385 1777 15419
rect 1777 15385 1811 15419
rect 1811 15385 1820 15419
rect 1768 15376 1820 15385
rect 4712 15376 4764 15428
rect 9036 15444 9088 15496
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 4436 15308 4488 15360
rect 5448 15308 5500 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 10232 15376 10284 15428
rect 11520 15444 11572 15496
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 12072 15419 12124 15428
rect 12072 15385 12081 15419
rect 12081 15385 12115 15419
rect 12115 15385 12124 15419
rect 12072 15376 12124 15385
rect 12532 15376 12584 15428
rect 7104 15308 7156 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 10324 15308 10376 15360
rect 10784 15308 10836 15360
rect 10968 15308 11020 15360
rect 11428 15308 11480 15360
rect 11796 15308 11848 15360
rect 14004 15308 14056 15360
rect 14096 15351 14148 15360
rect 14096 15317 14105 15351
rect 14105 15317 14139 15351
rect 14139 15317 14148 15351
rect 14096 15308 14148 15317
rect 3507 15206 3559 15258
rect 3571 15206 3623 15258
rect 3635 15206 3687 15258
rect 3699 15206 3751 15258
rect 3763 15206 3815 15258
rect 7302 15206 7354 15258
rect 7366 15206 7418 15258
rect 7430 15206 7482 15258
rect 7494 15206 7546 15258
rect 7558 15206 7610 15258
rect 11097 15206 11149 15258
rect 11161 15206 11213 15258
rect 11225 15206 11277 15258
rect 11289 15206 11341 15258
rect 11353 15206 11405 15258
rect 14892 15206 14944 15258
rect 14956 15206 15008 15258
rect 15020 15206 15072 15258
rect 15084 15206 15136 15258
rect 15148 15206 15200 15258
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 5264 15104 5316 15156
rect 5724 15104 5776 15156
rect 5448 15036 5500 15088
rect 7656 15104 7708 15156
rect 8944 15104 8996 15156
rect 9772 15104 9824 15156
rect 3976 14968 4028 15020
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 9956 15036 10008 15088
rect 11612 15104 11664 15156
rect 12532 15104 12584 15156
rect 14096 15104 14148 15156
rect 14648 15104 14700 15156
rect 13820 15036 13872 15088
rect 3884 14900 3936 14952
rect 7012 14900 7064 14952
rect 2688 14764 2740 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 13084 14968 13136 15020
rect 8484 14764 8536 14816
rect 9312 14764 9364 14816
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 14004 14968 14056 15020
rect 11428 14832 11480 14884
rect 12808 14764 12860 14816
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 2847 14662 2899 14714
rect 2911 14662 2963 14714
rect 2975 14662 3027 14714
rect 3039 14662 3091 14714
rect 3103 14662 3155 14714
rect 6642 14662 6694 14714
rect 6706 14662 6758 14714
rect 6770 14662 6822 14714
rect 6834 14662 6886 14714
rect 6898 14662 6950 14714
rect 10437 14662 10489 14714
rect 10501 14662 10553 14714
rect 10565 14662 10617 14714
rect 10629 14662 10681 14714
rect 10693 14662 10745 14714
rect 14232 14662 14284 14714
rect 14296 14662 14348 14714
rect 14360 14662 14412 14714
rect 14424 14662 14476 14714
rect 14488 14662 14540 14714
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 4252 14560 4304 14612
rect 5540 14560 5592 14612
rect 2780 14424 2832 14476
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 7012 14560 7064 14612
rect 8300 14560 8352 14612
rect 9864 14560 9916 14612
rect 10324 14492 10376 14544
rect 4528 14424 4580 14433
rect 6552 14424 6604 14476
rect 9312 14424 9364 14476
rect 10232 14424 10284 14476
rect 3884 14356 3936 14408
rect 4252 14356 4304 14408
rect 4436 14356 4488 14408
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 5816 14356 5868 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 11060 14356 11112 14408
rect 4344 14220 4396 14272
rect 5540 14220 5592 14272
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 5908 14288 5960 14340
rect 9220 14331 9272 14340
rect 9220 14297 9229 14331
rect 9229 14297 9263 14331
rect 9263 14297 9272 14331
rect 9220 14288 9272 14297
rect 9956 14288 10008 14340
rect 13820 14560 13872 14612
rect 11520 14356 11572 14408
rect 11888 14356 11940 14408
rect 12532 14356 12584 14408
rect 13636 14331 13688 14340
rect 13636 14297 13645 14331
rect 13645 14297 13679 14331
rect 13679 14297 13688 14331
rect 13636 14288 13688 14297
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 12164 14263 12216 14272
rect 12164 14229 12173 14263
rect 12173 14229 12207 14263
rect 12207 14229 12216 14263
rect 12164 14220 12216 14229
rect 3507 14118 3559 14170
rect 3571 14118 3623 14170
rect 3635 14118 3687 14170
rect 3699 14118 3751 14170
rect 3763 14118 3815 14170
rect 7302 14118 7354 14170
rect 7366 14118 7418 14170
rect 7430 14118 7482 14170
rect 7494 14118 7546 14170
rect 7558 14118 7610 14170
rect 11097 14118 11149 14170
rect 11161 14118 11213 14170
rect 11225 14118 11277 14170
rect 11289 14118 11341 14170
rect 11353 14118 11405 14170
rect 14892 14118 14944 14170
rect 14956 14118 15008 14170
rect 15020 14118 15072 14170
rect 15084 14118 15136 14170
rect 15148 14118 15200 14170
rect 2688 13948 2740 14000
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 5724 14016 5776 14068
rect 6460 14016 6512 14068
rect 7656 14016 7708 14068
rect 9036 14016 9088 14068
rect 9772 14016 9824 14068
rect 10784 14016 10836 14068
rect 11796 14016 11848 14068
rect 11888 14016 11940 14068
rect 12164 14016 12216 14068
rect 3884 13880 3936 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 6368 13948 6420 14000
rect 4804 13880 4856 13889
rect 8484 13880 8536 13932
rect 10324 13880 10376 13932
rect 12716 13991 12768 14000
rect 12716 13957 12725 13991
rect 12725 13957 12759 13991
rect 12759 13957 12768 13991
rect 12716 13948 12768 13957
rect 12808 13991 12860 14000
rect 12808 13957 12817 13991
rect 12817 13957 12851 13991
rect 12851 13957 12860 13991
rect 12808 13948 12860 13957
rect 5080 13812 5132 13864
rect 7012 13812 7064 13864
rect 5908 13744 5960 13796
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 12992 13812 13044 13864
rect 13636 14016 13688 14068
rect 9864 13744 9916 13796
rect 10048 13744 10100 13796
rect 12808 13744 12860 13796
rect 2780 13676 2832 13728
rect 3240 13676 3292 13728
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 2847 13574 2899 13626
rect 2911 13574 2963 13626
rect 2975 13574 3027 13626
rect 3039 13574 3091 13626
rect 3103 13574 3155 13626
rect 6642 13574 6694 13626
rect 6706 13574 6758 13626
rect 6770 13574 6822 13626
rect 6834 13574 6886 13626
rect 6898 13574 6950 13626
rect 10437 13574 10489 13626
rect 10501 13574 10553 13626
rect 10565 13574 10617 13626
rect 10629 13574 10681 13626
rect 10693 13574 10745 13626
rect 14232 13574 14284 13626
rect 14296 13574 14348 13626
rect 14360 13574 14412 13626
rect 14424 13574 14476 13626
rect 14488 13574 14540 13626
rect 2780 13472 2832 13524
rect 5080 13472 5132 13524
rect 12072 13472 12124 13524
rect 5540 13336 5592 13388
rect 13360 13472 13412 13524
rect 4344 13268 4396 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6644 13268 6696 13320
rect 12624 13336 12676 13388
rect 4252 13200 4304 13252
rect 4712 13132 4764 13184
rect 12716 13200 12768 13252
rect 5724 13132 5776 13184
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 3507 13030 3559 13082
rect 3571 13030 3623 13082
rect 3635 13030 3687 13082
rect 3699 13030 3751 13082
rect 3763 13030 3815 13082
rect 7302 13030 7354 13082
rect 7366 13030 7418 13082
rect 7430 13030 7482 13082
rect 7494 13030 7546 13082
rect 7558 13030 7610 13082
rect 11097 13030 11149 13082
rect 11161 13030 11213 13082
rect 11225 13030 11277 13082
rect 11289 13030 11341 13082
rect 11353 13030 11405 13082
rect 14892 13030 14944 13082
rect 14956 13030 15008 13082
rect 15020 13030 15072 13082
rect 15084 13030 15136 13082
rect 15148 13030 15200 13082
rect 6552 12928 6604 12980
rect 6644 12928 6696 12980
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 11888 12928 11940 12980
rect 12440 12928 12492 12980
rect 12532 12860 12584 12912
rect 5908 12792 5960 12844
rect 7564 12792 7616 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 3240 12724 3292 12776
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 7840 12724 7892 12776
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 2847 12486 2899 12538
rect 2911 12486 2963 12538
rect 2975 12486 3027 12538
rect 3039 12486 3091 12538
rect 3103 12486 3155 12538
rect 6642 12486 6694 12538
rect 6706 12486 6758 12538
rect 6770 12486 6822 12538
rect 6834 12486 6886 12538
rect 6898 12486 6950 12538
rect 10437 12486 10489 12538
rect 10501 12486 10553 12538
rect 10565 12486 10617 12538
rect 10629 12486 10681 12538
rect 10693 12486 10745 12538
rect 14232 12486 14284 12538
rect 14296 12486 14348 12538
rect 14360 12486 14412 12538
rect 14424 12486 14476 12538
rect 14488 12486 14540 12538
rect 4344 12384 4396 12436
rect 9864 12384 9916 12436
rect 1768 12248 1820 12300
rect 4712 12248 4764 12300
rect 5816 12291 5868 12300
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 6092 12248 6144 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 8024 12248 8076 12300
rect 12624 12248 12676 12300
rect 3332 12180 3384 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 7196 12180 7248 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 9680 12180 9732 12232
rect 13360 12180 13412 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 14740 12180 14792 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 2688 12044 2740 12096
rect 2964 12087 3016 12096
rect 2964 12053 2973 12087
rect 2973 12053 3007 12087
rect 3007 12053 3016 12087
rect 2964 12044 3016 12053
rect 7012 12044 7064 12096
rect 7380 12044 7432 12096
rect 8392 12044 8444 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11796 12044 11848 12096
rect 13544 12044 13596 12096
rect 14556 12044 14608 12096
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 3507 11942 3559 11994
rect 3571 11942 3623 11994
rect 3635 11942 3687 11994
rect 3699 11942 3751 11994
rect 3763 11942 3815 11994
rect 7302 11942 7354 11994
rect 7366 11942 7418 11994
rect 7430 11942 7482 11994
rect 7494 11942 7546 11994
rect 7558 11942 7610 11994
rect 11097 11942 11149 11994
rect 11161 11942 11213 11994
rect 11225 11942 11277 11994
rect 11289 11942 11341 11994
rect 11353 11942 11405 11994
rect 14892 11942 14944 11994
rect 14956 11942 15008 11994
rect 15020 11942 15072 11994
rect 15084 11942 15136 11994
rect 15148 11942 15200 11994
rect 1676 11840 1728 11892
rect 3424 11704 3476 11756
rect 7196 11840 7248 11892
rect 7196 11704 7248 11756
rect 10692 11840 10744 11892
rect 8484 11772 8536 11824
rect 9864 11772 9916 11824
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 9956 11704 10008 11756
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 6092 11568 6144 11620
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 9680 11500 9732 11552
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 14740 11704 14792 11756
rect 11520 11636 11572 11688
rect 12348 11636 12400 11688
rect 13544 11636 13596 11688
rect 15292 11772 15344 11824
rect 10324 11500 10376 11552
rect 10876 11500 10928 11552
rect 14648 11500 14700 11552
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 2847 11398 2899 11450
rect 2911 11398 2963 11450
rect 2975 11398 3027 11450
rect 3039 11398 3091 11450
rect 3103 11398 3155 11450
rect 6642 11398 6694 11450
rect 6706 11398 6758 11450
rect 6770 11398 6822 11450
rect 6834 11398 6886 11450
rect 6898 11398 6950 11450
rect 10437 11398 10489 11450
rect 10501 11398 10553 11450
rect 10565 11398 10617 11450
rect 10629 11398 10681 11450
rect 10693 11398 10745 11450
rect 14232 11398 14284 11450
rect 14296 11398 14348 11450
rect 14360 11398 14412 11450
rect 14424 11398 14476 11450
rect 14488 11398 14540 11450
rect 2780 11296 2832 11348
rect 3332 11296 3384 11348
rect 6460 11296 6512 11348
rect 7748 11296 7800 11348
rect 8208 11296 8260 11348
rect 8392 11296 8444 11348
rect 8576 11296 8628 11348
rect 10876 11296 10928 11348
rect 10968 11296 11020 11348
rect 6092 11160 6144 11212
rect 8300 11160 8352 11212
rect 9772 11160 9824 11212
rect 11520 11160 11572 11212
rect 12624 11296 12676 11348
rect 14556 11296 14608 11348
rect 15844 11339 15896 11348
rect 15844 11305 15853 11339
rect 15853 11305 15887 11339
rect 15887 11305 15896 11339
rect 15844 11296 15896 11305
rect 13820 11228 13872 11280
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 3148 11024 3200 11076
rect 6368 11024 6420 11076
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 11796 11092 11848 11144
rect 12532 11092 12584 11144
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 15384 11160 15436 11212
rect 9772 11024 9824 11076
rect 13728 11092 13780 11144
rect 2780 10999 2832 11008
rect 2780 10965 2789 10999
rect 2789 10965 2823 10999
rect 2823 10965 2832 10999
rect 2780 10956 2832 10965
rect 5908 10956 5960 11008
rect 8208 10956 8260 11008
rect 8484 10956 8536 11008
rect 9956 10956 10008 11008
rect 13912 11024 13964 11076
rect 11428 10956 11480 11008
rect 14740 10956 14792 11008
rect 3507 10854 3559 10906
rect 3571 10854 3623 10906
rect 3635 10854 3687 10906
rect 3699 10854 3751 10906
rect 3763 10854 3815 10906
rect 7302 10854 7354 10906
rect 7366 10854 7418 10906
rect 7430 10854 7482 10906
rect 7494 10854 7546 10906
rect 7558 10854 7610 10906
rect 11097 10854 11149 10906
rect 11161 10854 11213 10906
rect 11225 10854 11277 10906
rect 11289 10854 11341 10906
rect 11353 10854 11405 10906
rect 14892 10854 14944 10906
rect 14956 10854 15008 10906
rect 15020 10854 15072 10906
rect 15084 10854 15136 10906
rect 15148 10854 15200 10906
rect 3240 10752 3292 10804
rect 7196 10795 7248 10804
rect 7196 10761 7205 10795
rect 7205 10761 7239 10795
rect 7239 10761 7248 10795
rect 7196 10752 7248 10761
rect 3516 10684 3568 10736
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 4344 10616 4396 10668
rect 5908 10684 5960 10736
rect 9220 10684 9272 10736
rect 9772 10684 9824 10736
rect 10324 10684 10376 10736
rect 11428 10684 11480 10736
rect 6552 10480 6604 10532
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7196 10548 7248 10600
rect 8208 10616 8260 10668
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 9404 10616 9456 10668
rect 12348 10616 12400 10668
rect 13452 10616 13504 10668
rect 13728 10684 13780 10736
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 13820 10684 13872 10693
rect 14832 10616 14884 10668
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 7104 10412 7156 10464
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 10048 10412 10100 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 2847 10310 2899 10362
rect 2911 10310 2963 10362
rect 2975 10310 3027 10362
rect 3039 10310 3091 10362
rect 3103 10310 3155 10362
rect 6642 10310 6694 10362
rect 6706 10310 6758 10362
rect 6770 10310 6822 10362
rect 6834 10310 6886 10362
rect 6898 10310 6950 10362
rect 10437 10310 10489 10362
rect 10501 10310 10553 10362
rect 10565 10310 10617 10362
rect 10629 10310 10681 10362
rect 10693 10310 10745 10362
rect 14232 10310 14284 10362
rect 14296 10310 14348 10362
rect 14360 10310 14412 10362
rect 14424 10310 14476 10362
rect 14488 10310 14540 10362
rect 2504 10208 2556 10260
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 2320 10004 2372 10056
rect 3976 10208 4028 10260
rect 6092 10208 6144 10260
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 8300 10208 8352 10260
rect 8484 10140 8536 10192
rect 9220 10208 9272 10260
rect 9496 10208 9548 10260
rect 10140 10208 10192 10260
rect 12348 10208 12400 10260
rect 13912 10208 13964 10260
rect 15384 10208 15436 10260
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 3884 10047 3936 10056
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 7748 10072 7800 10124
rect 7656 10004 7708 10056
rect 9680 10072 9732 10124
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 14096 10140 14148 10192
rect 14556 10072 14608 10124
rect 8208 9936 8260 9988
rect 2780 9868 2832 9920
rect 6920 9868 6972 9920
rect 7104 9868 7156 9920
rect 7748 9868 7800 9920
rect 8116 9868 8168 9920
rect 9220 10004 9272 10056
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 10324 10004 10376 10056
rect 10968 10004 11020 10056
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 10600 9936 10652 9988
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 8760 9868 8812 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 3507 9766 3559 9818
rect 3571 9766 3623 9818
rect 3635 9766 3687 9818
rect 3699 9766 3751 9818
rect 3763 9766 3815 9818
rect 7302 9766 7354 9818
rect 7366 9766 7418 9818
rect 7430 9766 7482 9818
rect 7494 9766 7546 9818
rect 7558 9766 7610 9818
rect 11097 9766 11149 9818
rect 11161 9766 11213 9818
rect 11225 9766 11277 9818
rect 11289 9766 11341 9818
rect 11353 9766 11405 9818
rect 14892 9766 14944 9818
rect 14956 9766 15008 9818
rect 15020 9766 15072 9818
rect 15084 9766 15136 9818
rect 15148 9766 15200 9818
rect 2044 9664 2096 9716
rect 3792 9664 3844 9716
rect 4344 9664 4396 9716
rect 7104 9664 7156 9716
rect 7196 9664 7248 9716
rect 7656 9664 7708 9716
rect 3424 9596 3476 9648
rect 4528 9596 4580 9648
rect 6552 9596 6604 9648
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 4528 9460 4580 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 7196 9528 7248 9580
rect 3700 9324 3752 9376
rect 5816 9324 5868 9376
rect 6552 9324 6604 9376
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 8300 9596 8352 9648
rect 10324 9664 10376 9716
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 14096 9664 14148 9716
rect 15476 9664 15528 9716
rect 8392 9528 8444 9580
rect 8576 9528 8628 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9496 9528 9548 9580
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 8208 9460 8260 9512
rect 10140 9460 10192 9512
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 11796 9528 11848 9580
rect 13452 9503 13504 9512
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 8484 9392 8536 9444
rect 13820 9460 13872 9512
rect 14740 9460 14792 9512
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 8116 9324 8168 9376
rect 10968 9324 11020 9376
rect 11244 9324 11296 9376
rect 15292 9324 15344 9376
rect 2847 9222 2899 9274
rect 2911 9222 2963 9274
rect 2975 9222 3027 9274
rect 3039 9222 3091 9274
rect 3103 9222 3155 9274
rect 6642 9222 6694 9274
rect 6706 9222 6758 9274
rect 6770 9222 6822 9274
rect 6834 9222 6886 9274
rect 6898 9222 6950 9274
rect 10437 9222 10489 9274
rect 10501 9222 10553 9274
rect 10565 9222 10617 9274
rect 10629 9222 10681 9274
rect 10693 9222 10745 9274
rect 14232 9222 14284 9274
rect 14296 9222 14348 9274
rect 14360 9222 14412 9274
rect 14424 9222 14476 9274
rect 14488 9222 14540 9274
rect 2320 9120 2372 9172
rect 3700 9052 3752 9104
rect 5356 9120 5408 9172
rect 6828 9052 6880 9104
rect 5816 8984 5868 9036
rect 6736 8984 6788 9036
rect 8392 9120 8444 9172
rect 9220 9120 9272 9172
rect 8576 8984 8628 9036
rect 3332 8848 3384 8900
rect 7196 8916 7248 8968
rect 8116 8916 8168 8968
rect 6460 8848 6512 8900
rect 4528 8780 4580 8832
rect 7748 8891 7800 8900
rect 7748 8857 7757 8891
rect 7757 8857 7791 8891
rect 7791 8857 7800 8891
rect 7748 8848 7800 8857
rect 8668 8916 8720 8968
rect 9772 9120 9824 9172
rect 14556 9120 14608 9172
rect 9220 8780 9272 8832
rect 9588 8984 9640 9036
rect 9680 8984 9732 9036
rect 14188 8984 14240 9036
rect 15384 9052 15436 9104
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 10232 8916 10284 8968
rect 10692 8916 10744 8968
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 15660 8984 15712 9036
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 10784 8848 10836 8900
rect 11244 8891 11296 8900
rect 11244 8857 11253 8891
rect 11253 8857 11287 8891
rect 11287 8857 11296 8891
rect 11244 8848 11296 8857
rect 14280 8848 14332 8900
rect 10600 8780 10652 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 14740 8780 14792 8832
rect 3507 8678 3559 8730
rect 3571 8678 3623 8730
rect 3635 8678 3687 8730
rect 3699 8678 3751 8730
rect 3763 8678 3815 8730
rect 7302 8678 7354 8730
rect 7366 8678 7418 8730
rect 7430 8678 7482 8730
rect 7494 8678 7546 8730
rect 7558 8678 7610 8730
rect 11097 8678 11149 8730
rect 11161 8678 11213 8730
rect 11225 8678 11277 8730
rect 11289 8678 11341 8730
rect 11353 8678 11405 8730
rect 14892 8678 14944 8730
rect 14956 8678 15008 8730
rect 15020 8678 15072 8730
rect 15084 8678 15136 8730
rect 15148 8678 15200 8730
rect 6828 8576 6880 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8208 8576 8260 8628
rect 9312 8576 9364 8628
rect 10232 8576 10284 8628
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 10968 8619 11020 8628
rect 10968 8585 10995 8619
rect 10995 8585 11020 8619
rect 10968 8576 11020 8585
rect 7104 8508 7156 8560
rect 8484 8440 8536 8492
rect 10600 8508 10652 8560
rect 11428 8508 11480 8560
rect 10140 8440 10192 8492
rect 5264 8372 5316 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 7748 8304 7800 8356
rect 9220 8304 9272 8356
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12900 8576 12952 8628
rect 13452 8576 13504 8628
rect 14280 8576 14332 8628
rect 15292 8576 15344 8628
rect 15568 8576 15620 8628
rect 14004 8508 14056 8560
rect 12808 8372 12860 8424
rect 14188 8372 14240 8424
rect 13268 8304 13320 8356
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 10968 8279 11020 8288
rect 10968 8245 10977 8279
rect 10977 8245 11011 8279
rect 11011 8245 11020 8279
rect 10968 8236 11020 8245
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 12256 8236 12308 8288
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 15844 8304 15896 8356
rect 14648 8236 14700 8288
rect 15476 8236 15528 8288
rect 2847 8134 2899 8186
rect 2911 8134 2963 8186
rect 2975 8134 3027 8186
rect 3039 8134 3091 8186
rect 3103 8134 3155 8186
rect 6642 8134 6694 8186
rect 6706 8134 6758 8186
rect 6770 8134 6822 8186
rect 6834 8134 6886 8186
rect 6898 8134 6950 8186
rect 10437 8134 10489 8186
rect 10501 8134 10553 8186
rect 10565 8134 10617 8186
rect 10629 8134 10681 8186
rect 10693 8134 10745 8186
rect 14232 8134 14284 8186
rect 14296 8134 14348 8186
rect 14360 8134 14412 8186
rect 14424 8134 14476 8186
rect 14488 8134 14540 8186
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3976 7828 4028 7880
rect 8024 8032 8076 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9128 8032 9180 8084
rect 9496 8032 9548 8084
rect 9864 8032 9916 8084
rect 10692 8032 10744 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 13268 8032 13320 8084
rect 14096 8032 14148 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 8208 7828 8260 7880
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 15476 7828 15528 7880
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 4528 7692 4580 7744
rect 6920 7692 6972 7744
rect 9588 7760 9640 7812
rect 11520 7760 11572 7812
rect 9220 7735 9272 7744
rect 9220 7701 9245 7735
rect 9245 7701 9272 7735
rect 9220 7692 9272 7701
rect 9864 7692 9916 7744
rect 10692 7692 10744 7744
rect 13820 7692 13872 7744
rect 3507 7590 3559 7642
rect 3571 7590 3623 7642
rect 3635 7590 3687 7642
rect 3699 7590 3751 7642
rect 3763 7590 3815 7642
rect 7302 7590 7354 7642
rect 7366 7590 7418 7642
rect 7430 7590 7482 7642
rect 7494 7590 7546 7642
rect 7558 7590 7610 7642
rect 11097 7590 11149 7642
rect 11161 7590 11213 7642
rect 11225 7590 11277 7642
rect 11289 7590 11341 7642
rect 11353 7590 11405 7642
rect 14892 7590 14944 7642
rect 14956 7590 15008 7642
rect 15020 7590 15072 7642
rect 15084 7590 15136 7642
rect 15148 7590 15200 7642
rect 2412 7488 2464 7540
rect 3148 7488 3200 7540
rect 3976 7488 4028 7540
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 7748 7488 7800 7540
rect 3332 7420 3384 7472
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 3056 7284 3108 7336
rect 6000 7420 6052 7472
rect 8392 7488 8444 7540
rect 9404 7488 9456 7540
rect 9956 7488 10008 7540
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 12900 7488 12952 7540
rect 11244 7420 11296 7472
rect 14004 7488 14056 7540
rect 14740 7488 14792 7540
rect 15384 7488 15436 7540
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 7196 7284 7248 7336
rect 11980 7352 12032 7404
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 13912 7284 13964 7336
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 7012 7148 7064 7200
rect 9404 7148 9456 7200
rect 11152 7148 11204 7200
rect 14096 7148 14148 7200
rect 14648 7284 14700 7336
rect 15384 7284 15436 7336
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 2847 7046 2899 7098
rect 2911 7046 2963 7098
rect 2975 7046 3027 7098
rect 3039 7046 3091 7098
rect 3103 7046 3155 7098
rect 6642 7046 6694 7098
rect 6706 7046 6758 7098
rect 6770 7046 6822 7098
rect 6834 7046 6886 7098
rect 6898 7046 6950 7098
rect 10437 7046 10489 7098
rect 10501 7046 10553 7098
rect 10565 7046 10617 7098
rect 10629 7046 10681 7098
rect 10693 7046 10745 7098
rect 14232 7046 14284 7098
rect 14296 7046 14348 7098
rect 14360 7046 14412 7098
rect 14424 7046 14476 7098
rect 14488 7046 14540 7098
rect 1952 6944 2004 6996
rect 11244 6987 11296 6996
rect 11244 6953 11253 6987
rect 11253 6953 11287 6987
rect 11287 6953 11296 6987
rect 11244 6944 11296 6953
rect 13912 6944 13964 6996
rect 15476 6944 15528 6996
rect 3332 6808 3384 6860
rect 6552 6808 6604 6860
rect 9864 6808 9916 6860
rect 10876 6808 10928 6860
rect 11980 6808 12032 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 11152 6740 11204 6792
rect 7196 6672 7248 6724
rect 2044 6604 2096 6656
rect 3424 6604 3476 6656
rect 4436 6604 4488 6656
rect 6460 6604 6512 6656
rect 11704 6604 11756 6656
rect 15384 6740 15436 6792
rect 14648 6672 14700 6724
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 3507 6502 3559 6554
rect 3571 6502 3623 6554
rect 3635 6502 3687 6554
rect 3699 6502 3751 6554
rect 3763 6502 3815 6554
rect 7302 6502 7354 6554
rect 7366 6502 7418 6554
rect 7430 6502 7482 6554
rect 7494 6502 7546 6554
rect 7558 6502 7610 6554
rect 11097 6502 11149 6554
rect 11161 6502 11213 6554
rect 11225 6502 11277 6554
rect 11289 6502 11341 6554
rect 11353 6502 11405 6554
rect 14892 6502 14944 6554
rect 14956 6502 15008 6554
rect 15020 6502 15072 6554
rect 15084 6502 15136 6554
rect 15148 6502 15200 6554
rect 1676 6400 1728 6452
rect 3332 6400 3384 6452
rect 8944 6400 8996 6452
rect 10968 6400 11020 6452
rect 15660 6400 15712 6452
rect 9220 6332 9272 6384
rect 10140 6332 10192 6384
rect 11428 6332 11480 6384
rect 2044 6264 2096 6316
rect 3424 6264 3476 6316
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 6460 6196 6512 6248
rect 9864 6264 9916 6316
rect 9956 6264 10008 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 9680 6196 9732 6248
rect 9772 6128 9824 6180
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 10876 6060 10928 6112
rect 2847 5958 2899 6010
rect 2911 5958 2963 6010
rect 2975 5958 3027 6010
rect 3039 5958 3091 6010
rect 3103 5958 3155 6010
rect 6642 5958 6694 6010
rect 6706 5958 6758 6010
rect 6770 5958 6822 6010
rect 6834 5958 6886 6010
rect 6898 5958 6950 6010
rect 10437 5958 10489 6010
rect 10501 5958 10553 6010
rect 10565 5958 10617 6010
rect 10629 5958 10681 6010
rect 10693 5958 10745 6010
rect 14232 5958 14284 6010
rect 14296 5958 14348 6010
rect 14360 5958 14412 6010
rect 14424 5958 14476 6010
rect 14488 5958 14540 6010
rect 4712 5856 4764 5908
rect 6368 5856 6420 5908
rect 5816 5720 5868 5772
rect 6276 5720 6328 5772
rect 7196 5831 7248 5840
rect 7196 5797 7205 5831
rect 7205 5797 7239 5831
rect 7239 5797 7248 5831
rect 7196 5788 7248 5797
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 10140 5856 10192 5908
rect 11980 5856 12032 5908
rect 14740 5856 14792 5908
rect 15844 5856 15896 5908
rect 7196 5652 7248 5704
rect 9496 5652 9548 5704
rect 9763 5673 9815 5704
rect 9763 5652 9771 5673
rect 9771 5652 9805 5673
rect 9805 5652 9815 5673
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10324 5652 10376 5704
rect 10968 5652 11020 5704
rect 12072 5516 12124 5568
rect 3507 5414 3559 5466
rect 3571 5414 3623 5466
rect 3635 5414 3687 5466
rect 3699 5414 3751 5466
rect 3763 5414 3815 5466
rect 7302 5414 7354 5466
rect 7366 5414 7418 5466
rect 7430 5414 7482 5466
rect 7494 5414 7546 5466
rect 7558 5414 7610 5466
rect 11097 5414 11149 5466
rect 11161 5414 11213 5466
rect 11225 5414 11277 5466
rect 11289 5414 11341 5466
rect 11353 5414 11405 5466
rect 14892 5414 14944 5466
rect 14956 5414 15008 5466
rect 15020 5414 15072 5466
rect 15084 5414 15136 5466
rect 15148 5414 15200 5466
rect 5816 5355 5868 5364
rect 3240 5244 3292 5296
rect 2228 5176 2280 5228
rect 5816 5321 5825 5355
rect 5825 5321 5859 5355
rect 5859 5321 5868 5355
rect 5816 5312 5868 5321
rect 9036 5312 9088 5364
rect 9588 5355 9640 5364
rect 9588 5321 9597 5355
rect 9597 5321 9631 5355
rect 9631 5321 9640 5355
rect 9588 5312 9640 5321
rect 10048 5312 10100 5364
rect 5816 5176 5868 5228
rect 6736 5108 6788 5160
rect 5172 5040 5224 5092
rect 9956 5244 10008 5296
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 9588 5176 9640 5228
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 11336 5287 11388 5296
rect 11336 5253 11345 5287
rect 11345 5253 11379 5287
rect 11379 5253 11388 5287
rect 11336 5244 11388 5253
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 4160 4972 4212 5024
rect 5632 4972 5684 5024
rect 8668 4972 8720 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 9680 4972 9732 5024
rect 10140 5040 10192 5092
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 10968 5108 11020 5160
rect 11336 5108 11388 5160
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 10416 4972 10468 5024
rect 10784 4972 10836 5024
rect 11428 4972 11480 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 2847 4870 2899 4922
rect 2911 4870 2963 4922
rect 2975 4870 3027 4922
rect 3039 4870 3091 4922
rect 3103 4870 3155 4922
rect 6642 4870 6694 4922
rect 6706 4870 6758 4922
rect 6770 4870 6822 4922
rect 6834 4870 6886 4922
rect 6898 4870 6950 4922
rect 10437 4870 10489 4922
rect 10501 4870 10553 4922
rect 10565 4870 10617 4922
rect 10629 4870 10681 4922
rect 10693 4870 10745 4922
rect 14232 4870 14284 4922
rect 14296 4870 14348 4922
rect 14360 4870 14412 4922
rect 14424 4870 14476 4922
rect 14488 4870 14540 4922
rect 3332 4768 3384 4820
rect 4436 4768 4488 4820
rect 6552 4768 6604 4820
rect 2688 4700 2740 4752
rect 4252 4564 4304 4616
rect 3240 4496 3292 4548
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 5632 4632 5684 4684
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 5172 4564 5224 4616
rect 7196 4768 7248 4820
rect 8668 4811 8720 4820
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 10968 4768 11020 4820
rect 11428 4768 11480 4820
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 11980 4632 12032 4684
rect 1952 4428 2004 4480
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 4344 4428 4396 4480
rect 6000 4496 6052 4548
rect 8208 4496 8260 4548
rect 5724 4428 5776 4480
rect 8116 4428 8168 4480
rect 9220 4428 9272 4480
rect 9864 4496 9916 4548
rect 10784 4496 10836 4548
rect 9588 4428 9640 4480
rect 11336 4428 11388 4480
rect 12900 4564 12952 4616
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 3507 4326 3559 4378
rect 3571 4326 3623 4378
rect 3635 4326 3687 4378
rect 3699 4326 3751 4378
rect 3763 4326 3815 4378
rect 7302 4326 7354 4378
rect 7366 4326 7418 4378
rect 7430 4326 7482 4378
rect 7494 4326 7546 4378
rect 7558 4326 7610 4378
rect 11097 4326 11149 4378
rect 11161 4326 11213 4378
rect 11225 4326 11277 4378
rect 11289 4326 11341 4378
rect 11353 4326 11405 4378
rect 14892 4326 14944 4378
rect 14956 4326 15008 4378
rect 15020 4326 15072 4378
rect 15084 4326 15136 4378
rect 15148 4326 15200 4378
rect 3240 4224 3292 4276
rect 9036 4267 9088 4276
rect 9036 4233 9045 4267
rect 9045 4233 9079 4267
rect 9079 4233 9088 4267
rect 9036 4224 9088 4233
rect 9128 4224 9180 4276
rect 9864 4224 9916 4276
rect 10784 4224 10836 4276
rect 2228 4156 2280 4208
rect 2320 4199 2372 4208
rect 2320 4165 2329 4199
rect 2329 4165 2363 4199
rect 2363 4165 2372 4199
rect 2320 4156 2372 4165
rect 3332 4156 3384 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2688 4020 2740 4072
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 5724 4088 5776 4140
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 4252 4020 4304 4072
rect 3056 3884 3108 3936
rect 3976 3884 4028 3936
rect 6092 4020 6144 4072
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 12900 4156 12952 4208
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 5908 3884 5960 3936
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 9680 4088 9732 4140
rect 11980 4088 12032 4140
rect 9496 4020 9548 4072
rect 11060 4020 11112 4072
rect 12808 4020 12860 4072
rect 9772 3884 9824 3936
rect 11428 3952 11480 4004
rect 12624 3884 12676 3936
rect 2847 3782 2899 3834
rect 2911 3782 2963 3834
rect 2975 3782 3027 3834
rect 3039 3782 3091 3834
rect 3103 3782 3155 3834
rect 6642 3782 6694 3834
rect 6706 3782 6758 3834
rect 6770 3782 6822 3834
rect 6834 3782 6886 3834
rect 6898 3782 6950 3834
rect 10437 3782 10489 3834
rect 10501 3782 10553 3834
rect 10565 3782 10617 3834
rect 10629 3782 10681 3834
rect 10693 3782 10745 3834
rect 14232 3782 14284 3834
rect 14296 3782 14348 3834
rect 14360 3782 14412 3834
rect 14424 3782 14476 3834
rect 14488 3782 14540 3834
rect 2228 3680 2280 3732
rect 4344 3680 4396 3732
rect 2044 3544 2096 3596
rect 5908 3680 5960 3732
rect 6092 3680 6144 3732
rect 7196 3680 7248 3732
rect 8668 3680 8720 3732
rect 10140 3680 10192 3732
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 12624 3680 12676 3732
rect 3332 3476 3384 3528
rect 3976 3476 4028 3528
rect 4252 3476 4304 3528
rect 5264 3476 5316 3528
rect 1952 3408 2004 3460
rect 5724 3408 5776 3460
rect 8116 3476 8168 3528
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 6000 3408 6052 3460
rect 9128 3544 9180 3596
rect 9588 3544 9640 3596
rect 10048 3544 10100 3596
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 12716 3476 12768 3528
rect 13820 3476 13872 3528
rect 9588 3408 9640 3460
rect 6736 3340 6788 3392
rect 9864 3340 9916 3392
rect 3507 3238 3559 3290
rect 3571 3238 3623 3290
rect 3635 3238 3687 3290
rect 3699 3238 3751 3290
rect 3763 3238 3815 3290
rect 7302 3238 7354 3290
rect 7366 3238 7418 3290
rect 7430 3238 7482 3290
rect 7494 3238 7546 3290
rect 7558 3238 7610 3290
rect 11097 3238 11149 3290
rect 11161 3238 11213 3290
rect 11225 3238 11277 3290
rect 11289 3238 11341 3290
rect 11353 3238 11405 3290
rect 14892 3238 14944 3290
rect 14956 3238 15008 3290
rect 15020 3238 15072 3290
rect 15084 3238 15136 3290
rect 15148 3238 15200 3290
rect 5816 3136 5868 3188
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 9680 3136 9732 3188
rect 9864 3136 9916 3188
rect 10968 3136 11020 3188
rect 11428 3136 11480 3188
rect 6736 3068 6788 3120
rect 5724 3000 5776 3052
rect 8208 3000 8260 3052
rect 10876 3000 10928 3052
rect 12624 3000 12676 3052
rect 13820 2932 13872 2984
rect 2847 2694 2899 2746
rect 2911 2694 2963 2746
rect 2975 2694 3027 2746
rect 3039 2694 3091 2746
rect 3103 2694 3155 2746
rect 6642 2694 6694 2746
rect 6706 2694 6758 2746
rect 6770 2694 6822 2746
rect 6834 2694 6886 2746
rect 6898 2694 6950 2746
rect 10437 2694 10489 2746
rect 10501 2694 10553 2746
rect 10565 2694 10617 2746
rect 10629 2694 10681 2746
rect 10693 2694 10745 2746
rect 14232 2694 14284 2746
rect 14296 2694 14348 2746
rect 14360 2694 14412 2746
rect 14424 2694 14476 2746
rect 14488 2694 14540 2746
rect 4436 2592 4488 2644
rect 13820 2456 13872 2508
rect 20 2388 72 2440
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 3507 2150 3559 2202
rect 3571 2150 3623 2202
rect 3635 2150 3687 2202
rect 3699 2150 3751 2202
rect 3763 2150 3815 2202
rect 7302 2150 7354 2202
rect 7366 2150 7418 2202
rect 7430 2150 7482 2202
rect 7494 2150 7546 2202
rect 7558 2150 7610 2202
rect 11097 2150 11149 2202
rect 11161 2150 11213 2202
rect 11225 2150 11277 2202
rect 11289 2150 11341 2202
rect 11353 2150 11405 2202
rect 14892 2150 14944 2202
rect 14956 2150 15008 2202
rect 15020 2150 15072 2202
rect 15084 2150 15136 2202
rect 15148 2150 15200 2202
<< metal2 >>
rect 9678 18774 9734 19574
rect 2847 16892 3155 16901
rect 2847 16890 2853 16892
rect 2909 16890 2933 16892
rect 2989 16890 3013 16892
rect 3069 16890 3093 16892
rect 3149 16890 3155 16892
rect 2909 16838 2911 16890
rect 3091 16838 3093 16890
rect 2847 16836 2853 16838
rect 2909 16836 2933 16838
rect 2989 16836 3013 16838
rect 3069 16836 3093 16838
rect 3149 16836 3155 16838
rect 2847 16827 3155 16836
rect 6642 16892 6950 16901
rect 6642 16890 6648 16892
rect 6704 16890 6728 16892
rect 6784 16890 6808 16892
rect 6864 16890 6888 16892
rect 6944 16890 6950 16892
rect 6704 16838 6706 16890
rect 6886 16838 6888 16890
rect 6642 16836 6648 16838
rect 6704 16836 6728 16838
rect 6784 16836 6808 16838
rect 6864 16836 6888 16838
rect 6944 16836 6950 16838
rect 6642 16827 6950 16836
rect 9692 16574 9720 18774
rect 10437 16892 10745 16901
rect 10437 16890 10443 16892
rect 10499 16890 10523 16892
rect 10579 16890 10603 16892
rect 10659 16890 10683 16892
rect 10739 16890 10745 16892
rect 10499 16838 10501 16890
rect 10681 16838 10683 16890
rect 10437 16836 10443 16838
rect 10499 16836 10523 16838
rect 10579 16836 10603 16838
rect 10659 16836 10683 16838
rect 10739 16836 10745 16838
rect 10437 16827 10745 16836
rect 14232 16892 14540 16901
rect 14232 16890 14238 16892
rect 14294 16890 14318 16892
rect 14374 16890 14398 16892
rect 14454 16890 14478 16892
rect 14534 16890 14540 16892
rect 14294 16838 14296 16890
rect 14476 16838 14478 16890
rect 14232 16836 14238 16838
rect 14294 16836 14318 16838
rect 14374 16836 14398 16838
rect 14454 16836 14478 16838
rect 14534 16836 14540 16838
rect 14232 16827 14540 16836
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 9864 16584 9916 16590
rect 9692 16546 9864 16574
rect 9864 16526 9916 16532
rect 3507 16348 3815 16357
rect 3507 16346 3513 16348
rect 3569 16346 3593 16348
rect 3649 16346 3673 16348
rect 3729 16346 3753 16348
rect 3809 16346 3815 16348
rect 3569 16294 3571 16346
rect 3751 16294 3753 16346
rect 3507 16292 3513 16294
rect 3569 16292 3593 16294
rect 3649 16292 3673 16294
rect 3729 16292 3753 16294
rect 3809 16292 3815 16294
rect 3507 16283 3815 16292
rect 7302 16348 7610 16357
rect 7302 16346 7308 16348
rect 7364 16346 7388 16348
rect 7444 16346 7468 16348
rect 7524 16346 7548 16348
rect 7604 16346 7610 16348
rect 7364 16294 7366 16346
rect 7546 16294 7548 16346
rect 7302 16292 7308 16294
rect 7364 16292 7388 16294
rect 7444 16292 7468 16294
rect 7524 16292 7548 16294
rect 7604 16292 7610 16294
rect 7302 16283 7610 16292
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 2847 15804 3155 15813
rect 2847 15802 2853 15804
rect 2909 15802 2933 15804
rect 2989 15802 3013 15804
rect 3069 15802 3093 15804
rect 3149 15802 3155 15804
rect 2909 15750 2911 15802
rect 3091 15750 3093 15802
rect 2847 15748 2853 15750
rect 2909 15748 2933 15750
rect 2989 15748 3013 15750
rect 3069 15748 3093 15750
rect 3149 15748 3155 15750
rect 2847 15739 3155 15748
rect 3988 15502 4016 15846
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1780 12306 1808 15370
rect 3507 15260 3815 15269
rect 3507 15258 3513 15260
rect 3569 15258 3593 15260
rect 3649 15258 3673 15260
rect 3729 15258 3753 15260
rect 3809 15258 3815 15260
rect 3569 15206 3571 15258
rect 3751 15206 3753 15258
rect 3507 15204 3513 15206
rect 3569 15204 3593 15206
rect 3649 15204 3673 15206
rect 3729 15204 3753 15206
rect 3809 15204 3815 15206
rect 3507 15195 3815 15204
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2700 14634 2728 14758
rect 2847 14716 3155 14725
rect 2847 14714 2853 14716
rect 2909 14714 2933 14716
rect 2989 14714 3013 14716
rect 3069 14714 3093 14716
rect 3149 14714 3155 14716
rect 2909 14662 2911 14714
rect 3091 14662 3093 14714
rect 2847 14660 2853 14662
rect 2909 14660 2933 14662
rect 2989 14660 3013 14662
rect 3069 14660 3093 14662
rect 3149 14660 3155 14662
rect 2847 14651 3155 14660
rect 2700 14606 2820 14634
rect 3896 14618 3924 14894
rect 2792 14482 2820 14606
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2700 13546 2728 13942
rect 2792 13734 2820 14418
rect 3884 14408 3936 14414
rect 3988 14396 4016 14962
rect 4264 14618 4292 15438
rect 4356 15162 4384 15982
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3936 14368 4016 14396
rect 4252 14408 4304 14414
rect 3884 14350 3936 14356
rect 4252 14350 4304 14356
rect 3507 14172 3815 14181
rect 3507 14170 3513 14172
rect 3569 14170 3593 14172
rect 3649 14170 3673 14172
rect 3729 14170 3753 14172
rect 3809 14170 3815 14172
rect 3569 14118 3571 14170
rect 3751 14118 3753 14170
rect 3507 14116 3513 14118
rect 3569 14116 3593 14118
rect 3649 14116 3673 14118
rect 3729 14116 3753 14118
rect 3809 14116 3815 14118
rect 3507 14107 3815 14116
rect 3896 13938 3924 14350
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 2847 13628 3155 13637
rect 2847 13626 2853 13628
rect 2909 13626 2933 13628
rect 2989 13626 3013 13628
rect 3069 13626 3093 13628
rect 3149 13626 3155 13628
rect 2909 13574 2911 13626
rect 3091 13574 3093 13626
rect 2847 13572 2853 13574
rect 2909 13572 2933 13574
rect 2989 13572 3013 13574
rect 3069 13572 3093 13574
rect 3149 13572 3155 13574
rect 2847 13563 3155 13572
rect 2700 13530 2820 13546
rect 2700 13524 2832 13530
rect 2700 13518 2780 13524
rect 2780 13466 2832 13472
rect 3252 12782 3280 13670
rect 4264 13258 4292 14350
rect 4356 14278 4384 15098
rect 4448 14414 4476 15302
rect 4540 14482 4568 15506
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4724 14074 4752 15370
rect 4816 14414 4844 15846
rect 5276 15162 5304 15982
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15706 6224 15846
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5460 15094 5488 15302
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5552 14618 5580 15438
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15162 5764 15302
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 6196 15026 6224 15506
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 6196 14414 6224 14962
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 13326 4384 13670
rect 4816 13326 4844 13874
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13530 5120 13806
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5552 13394 5580 14214
rect 5736 14074 5764 14214
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 3507 13084 3815 13093
rect 3507 13082 3513 13084
rect 3569 13082 3593 13084
rect 3649 13082 3673 13084
rect 3729 13082 3753 13084
rect 3809 13082 3815 13084
rect 3569 13030 3571 13082
rect 3751 13030 3753 13082
rect 3507 13028 3513 13030
rect 3569 13028 3593 13030
rect 3649 13028 3673 13030
rect 3729 13028 3753 13030
rect 3809 13028 3815 13030
rect 3507 13019 3815 13028
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 2847 12540 3155 12549
rect 2847 12538 2853 12540
rect 2909 12538 2933 12540
rect 2989 12538 3013 12540
rect 3069 12538 3093 12540
rect 3149 12538 3155 12540
rect 2909 12486 2911 12538
rect 3091 12486 3093 12538
rect 2847 12484 2853 12486
rect 2909 12484 2933 12486
rect 2989 12484 3013 12486
rect 3069 12484 3093 12486
rect 3149 12484 3155 12486
rect 2847 12475 3155 12484
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1780 11914 1808 12242
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 1688 11898 1808 11914
rect 1676 11892 1808 11898
rect 1728 11886 1808 11892
rect 1676 11834 1728 11840
rect 2700 11336 2728 12038
rect 2976 11694 3004 12038
rect 3252 11694 3280 12718
rect 4356 12442 4384 12718
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4724 12306 4752 13126
rect 5736 12434 5764 13126
rect 5552 12406 5764 12434
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 5552 12238 5580 12406
rect 5828 12306 5856 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 13802 5948 14282
rect 6380 14006 6408 15982
rect 6472 14074 6500 16050
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 6642 15804 6950 15813
rect 6642 15802 6648 15804
rect 6704 15802 6728 15804
rect 6784 15802 6808 15804
rect 6864 15802 6888 15804
rect 6944 15802 6950 15804
rect 6704 15750 6706 15802
rect 6886 15750 6888 15802
rect 6642 15748 6648 15750
rect 6704 15748 6728 15750
rect 6784 15748 6808 15750
rect 6864 15748 6888 15750
rect 6944 15748 6950 15750
rect 6642 15739 6950 15748
rect 7392 15706 7420 15982
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 15706 9076 15846
rect 9600 15706 9628 15982
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14482 6592 14758
rect 6642 14716 6950 14725
rect 6642 14714 6648 14716
rect 6704 14714 6728 14716
rect 6784 14714 6808 14716
rect 6864 14714 6888 14716
rect 6944 14714 6950 14716
rect 6704 14662 6706 14714
rect 6886 14662 6888 14714
rect 6642 14660 6648 14662
rect 6704 14660 6728 14662
rect 6784 14660 6808 14662
rect 6864 14660 6888 14662
rect 6944 14660 6950 14662
rect 6642 14651 6950 14660
rect 7024 14618 7052 14894
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 7024 13870 7052 14554
rect 7116 14464 7144 15302
rect 7302 15260 7610 15269
rect 7302 15258 7308 15260
rect 7364 15258 7388 15260
rect 7444 15258 7468 15260
rect 7524 15258 7548 15260
rect 7604 15258 7610 15260
rect 7364 15206 7366 15258
rect 7546 15206 7548 15258
rect 7302 15204 7308 15206
rect 7364 15204 7388 15206
rect 7444 15204 7468 15206
rect 7524 15204 7548 15206
rect 7604 15204 7610 15206
rect 7302 15195 7610 15204
rect 7668 15162 7696 15302
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7116 14436 7236 14464
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 12850 5948 13738
rect 6642 13628 6950 13637
rect 6642 13626 6648 13628
rect 6704 13626 6728 13628
rect 6784 13626 6808 13628
rect 6864 13626 6888 13628
rect 6944 13626 6950 13628
rect 6704 13574 6706 13626
rect 6886 13574 6888 13626
rect 6642 13572 6648 13574
rect 6704 13572 6728 13574
rect 6784 13572 6808 13574
rect 6864 13572 6888 13574
rect 6944 13572 6950 13574
rect 6642 13563 6950 13572
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6564 12986 6592 13262
rect 6656 12986 6684 13262
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12986 6776 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 2847 11452 3155 11461
rect 2847 11450 2853 11452
rect 2909 11450 2933 11452
rect 2989 11450 3013 11452
rect 3069 11450 3093 11452
rect 3149 11450 3155 11452
rect 2909 11398 2911 11450
rect 3091 11398 3093 11450
rect 2847 11396 2853 11398
rect 2909 11396 2933 11398
rect 2989 11396 3013 11398
rect 3069 11396 3093 11398
rect 3149 11396 3155 11398
rect 2847 11387 3155 11396
rect 2780 11348 2832 11354
rect 2700 11308 2780 11336
rect 2780 11290 2832 11296
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 10266 2544 10542
rect 2792 10418 2820 10950
rect 3160 10554 3188 11018
rect 3252 10810 3280 11630
rect 3344 11354 3372 12174
rect 3507 11996 3815 12005
rect 3507 11994 3513 11996
rect 3569 11994 3593 11996
rect 3649 11994 3673 11996
rect 3729 11994 3753 11996
rect 3809 11994 3815 11996
rect 3569 11942 3571 11994
rect 3751 11942 3753 11994
rect 3507 11940 3513 11942
rect 3569 11940 3593 11942
rect 3649 11940 3673 11942
rect 3729 11940 3753 11942
rect 3809 11940 3815 11942
rect 3507 11931 3815 11940
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3436 10724 3464 11698
rect 5920 11014 5948 12786
rect 7024 12782 7052 13806
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6642 12540 6950 12549
rect 6642 12538 6648 12540
rect 6704 12538 6728 12540
rect 6784 12538 6808 12540
rect 6864 12538 6888 12540
rect 6944 12538 6950 12540
rect 6704 12486 6706 12538
rect 6886 12486 6888 12538
rect 6642 12484 6648 12486
rect 6704 12484 6728 12486
rect 6784 12484 6808 12486
rect 6864 12484 6888 12486
rect 6944 12484 6950 12486
rect 6642 12475 6950 12484
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6104 11626 6132 12242
rect 7208 12238 7236 14436
rect 7302 14172 7610 14181
rect 7302 14170 7308 14172
rect 7364 14170 7388 14172
rect 7444 14170 7468 14172
rect 7524 14170 7548 14172
rect 7604 14170 7610 14172
rect 7364 14118 7366 14170
rect 7546 14118 7548 14170
rect 7302 14116 7308 14118
rect 7364 14116 7388 14118
rect 7444 14116 7468 14118
rect 7524 14116 7548 14118
rect 7604 14116 7610 14118
rect 7302 14107 7610 14116
rect 7668 14074 7696 15098
rect 8312 14618 8340 15438
rect 8496 14822 8524 15438
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15162 8984 15302
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 8496 13938 8524 14758
rect 9048 14074 9076 15438
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9232 14346 9260 15302
rect 9784 15162 9812 15982
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15502 9904 15846
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9876 15042 9904 15438
rect 9784 15014 9904 15042
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14482 9352 14758
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9784 14074 9812 15014
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14618 9904 14894
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9968 14346 9996 15030
rect 10060 14464 10088 15506
rect 10244 15434 10272 16594
rect 11097 16348 11405 16357
rect 11097 16346 11103 16348
rect 11159 16346 11183 16348
rect 11239 16346 11263 16348
rect 11319 16346 11343 16348
rect 11399 16346 11405 16348
rect 11159 16294 11161 16346
rect 11341 16294 11343 16346
rect 11097 16292 11103 16294
rect 11159 16292 11183 16294
rect 11239 16292 11263 16294
rect 11319 16292 11343 16294
rect 11399 16292 11405 16294
rect 11097 16283 11405 16292
rect 14892 16348 15200 16357
rect 14892 16346 14898 16348
rect 14954 16346 14978 16348
rect 15034 16346 15058 16348
rect 15114 16346 15138 16348
rect 15194 16346 15200 16348
rect 14954 16294 14956 16346
rect 15136 16294 15138 16346
rect 14892 16292 14898 16294
rect 14954 16292 14978 16294
rect 15034 16292 15058 16294
rect 15114 16292 15138 16294
rect 15194 16292 15200 16294
rect 14892 16283 15200 16292
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 10437 15804 10745 15813
rect 10437 15802 10443 15804
rect 10499 15802 10523 15804
rect 10579 15802 10603 15804
rect 10659 15802 10683 15804
rect 10739 15802 10745 15804
rect 10499 15750 10501 15802
rect 10681 15750 10683 15802
rect 10437 15748 10443 15750
rect 10499 15748 10523 15750
rect 10579 15748 10603 15750
rect 10659 15748 10683 15750
rect 10739 15748 10745 15750
rect 10437 15739 10745 15748
rect 11532 15638 11560 15846
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 10336 14550 10364 15302
rect 10437 14716 10745 14725
rect 10437 14714 10443 14716
rect 10499 14714 10523 14716
rect 10579 14714 10603 14716
rect 10659 14714 10683 14716
rect 10739 14714 10745 14716
rect 10499 14662 10501 14714
rect 10681 14662 10683 14714
rect 10437 14660 10443 14662
rect 10499 14660 10523 14662
rect 10579 14660 10603 14662
rect 10659 14660 10683 14662
rect 10739 14660 10745 14662
rect 10437 14651 10745 14660
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10232 14476 10284 14482
rect 10060 14436 10232 14464
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 7302 13084 7610 13093
rect 7302 13082 7308 13084
rect 7364 13082 7388 13084
rect 7444 13082 7468 13084
rect 7524 13082 7548 13084
rect 7604 13082 7610 13084
rect 7364 13030 7366 13082
rect 7546 13030 7548 13082
rect 7302 13028 7308 13030
rect 7364 13028 7388 13030
rect 7444 13028 7468 13030
rect 7524 13028 7548 13030
rect 7604 13028 7610 13030
rect 7302 13019 7610 13028
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12306 7604 12786
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7852 12434 7880 12718
rect 7668 12406 7880 12434
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7012 12096 7064 12102
rect 7380 12096 7432 12102
rect 7012 12038 7064 12044
rect 7208 12056 7380 12084
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6104 11218 6132 11562
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11354 6500 11494
rect 6642 11452 6950 11461
rect 6642 11450 6648 11452
rect 6704 11450 6728 11452
rect 6784 11450 6808 11452
rect 6864 11450 6888 11452
rect 6944 11450 6950 11452
rect 6704 11398 6706 11450
rect 6886 11398 6888 11450
rect 6642 11396 6648 11398
rect 6704 11396 6728 11398
rect 6784 11396 6808 11398
rect 6864 11396 6888 11398
rect 6944 11396 6950 11398
rect 6642 11387 6950 11396
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 3507 10908 3815 10917
rect 3507 10906 3513 10908
rect 3569 10906 3593 10908
rect 3649 10906 3673 10908
rect 3729 10906 3753 10908
rect 3809 10906 3815 10908
rect 3569 10854 3571 10906
rect 3751 10854 3753 10906
rect 3507 10852 3513 10854
rect 3569 10852 3593 10854
rect 3649 10852 3673 10854
rect 3729 10852 3753 10854
rect 3809 10852 3815 10854
rect 3507 10843 3815 10852
rect 5920 10742 5948 10950
rect 3516 10736 3568 10742
rect 3436 10696 3516 10724
rect 3160 10526 3280 10554
rect 2700 10390 2820 10418
rect 2700 10282 2728 10390
rect 2847 10364 3155 10373
rect 2847 10362 2853 10364
rect 2909 10362 2933 10364
rect 2989 10362 3013 10364
rect 3069 10362 3093 10364
rect 3149 10362 3155 10364
rect 2909 10310 2911 10362
rect 3091 10310 3093 10362
rect 2847 10308 2853 10310
rect 2909 10308 2933 10310
rect 2989 10308 3013 10310
rect 3069 10308 3093 10310
rect 3149 10308 3155 10310
rect 2847 10299 3155 10308
rect 2504 10260 2556 10266
rect 2700 10254 2820 10282
rect 2504 10202 2556 10208
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2056 9722 2084 9998
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2332 9178 2360 9998
rect 2792 9926 2820 10254
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2847 9276 3155 9285
rect 2847 9274 2853 9276
rect 2909 9274 2933 9276
rect 2989 9274 3013 9276
rect 3069 9274 3093 9276
rect 3149 9274 3155 9276
rect 2909 9222 2911 9274
rect 3091 9222 3093 9274
rect 2847 9220 2853 9222
rect 2909 9220 2933 9222
rect 2989 9220 3013 9222
rect 3069 9220 3093 9222
rect 3149 9220 3155 9222
rect 2847 9211 3155 9220
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2847 8188 3155 8197
rect 2847 8186 2853 8188
rect 2909 8186 2933 8188
rect 2989 8186 3013 8188
rect 3069 8186 3093 8188
rect 3149 8186 3155 8188
rect 2909 8134 2911 8186
rect 3091 8134 3093 8186
rect 2847 8132 2853 8134
rect 2909 8132 2933 8134
rect 2989 8132 3013 8134
rect 3069 8132 3093 8134
rect 3149 8132 3155 8134
rect 2847 8123 3155 8132
rect 3252 7954 3280 10526
rect 3436 9654 3464 10696
rect 3516 10678 3568 10684
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10266 4016 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3507 9820 3815 9829
rect 3507 9818 3513 9820
rect 3569 9818 3593 9820
rect 3649 9818 3673 9820
rect 3729 9818 3753 9820
rect 3809 9818 3815 9820
rect 3569 9766 3571 9818
rect 3751 9766 3753 9818
rect 3507 9764 3513 9766
rect 3569 9764 3593 9766
rect 3649 9764 3673 9766
rect 3729 9764 3753 9766
rect 3809 9764 3815 9766
rect 3507 9755 3815 9764
rect 3792 9716 3844 9722
rect 3896 9704 3924 9998
rect 4356 9722 4384 10610
rect 6104 10266 6132 11154
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 3844 9676 3924 9704
rect 4344 9716 4396 9722
rect 3792 9658 3844 9664
rect 4344 9658 4396 9664
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 9110 3740 9318
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2424 7546 2452 7686
rect 3160 7546 3188 7686
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3252 7426 3280 7890
rect 3344 7478 3372 8842
rect 3507 8732 3815 8741
rect 3507 8730 3513 8732
rect 3569 8730 3593 8732
rect 3649 8730 3673 8732
rect 3729 8730 3753 8732
rect 3809 8730 3815 8732
rect 3569 8678 3571 8730
rect 3751 8678 3753 8730
rect 3507 8676 3513 8678
rect 3569 8676 3593 8678
rect 3649 8676 3673 8678
rect 3729 8676 3753 8678
rect 3809 8676 3815 8678
rect 3507 8667 3815 8676
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3507 7644 3815 7653
rect 3507 7642 3513 7644
rect 3569 7642 3593 7644
rect 3649 7642 3673 7644
rect 3729 7642 3753 7644
rect 3809 7642 3815 7644
rect 3569 7590 3571 7642
rect 3751 7590 3753 7642
rect 3507 7588 3513 7590
rect 3569 7588 3593 7590
rect 3649 7588 3673 7590
rect 3729 7588 3753 7590
rect 3809 7588 3815 7590
rect 3507 7579 3815 7588
rect 3988 7546 4016 7822
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3068 7398 3280 7426
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3068 7342 3096 7398
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 1688 6458 1716 7278
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 7002 1992 7142
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2056 6662 2084 7278
rect 2847 7100 3155 7109
rect 2847 7098 2853 7100
rect 2909 7098 2933 7100
rect 2989 7098 3013 7100
rect 3069 7098 3093 7100
rect 3149 7098 3155 7100
rect 2909 7046 2911 7098
rect 3091 7046 3093 7098
rect 2847 7044 2853 7046
rect 2909 7044 2933 7046
rect 2989 7044 3013 7046
rect 3069 7044 3093 7046
rect 3149 7044 3155 7046
rect 2847 7035 3155 7044
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2056 6322 2084 6598
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 3466 1992 4422
rect 2056 4146 2084 6258
rect 2847 6012 3155 6021
rect 2847 6010 2853 6012
rect 2909 6010 2933 6012
rect 2989 6010 3013 6012
rect 3069 6010 3093 6012
rect 3149 6010 3155 6012
rect 2909 5958 2911 6010
rect 3091 5958 3093 6010
rect 2847 5956 2853 5958
rect 2909 5956 2933 5958
rect 2989 5956 3013 5958
rect 3069 5956 3093 5958
rect 3149 5956 3155 5958
rect 2847 5947 3155 5956
rect 3252 5302 3280 7398
rect 3344 6866 3372 7414
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 6458 3372 6802
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2240 4214 2268 5170
rect 2847 4924 3155 4933
rect 2847 4922 2853 4924
rect 2909 4922 2933 4924
rect 2989 4922 3013 4924
rect 3069 4922 3093 4924
rect 3149 4922 3155 4924
rect 2909 4870 2911 4922
rect 3091 4870 3093 4922
rect 2847 4868 2853 4870
rect 2909 4868 2933 4870
rect 2989 4868 3013 4870
rect 3069 4868 3093 4870
rect 3149 4868 3155 4870
rect 2847 4859 3155 4868
rect 2688 4752 2740 4758
rect 3252 4706 3280 5238
rect 3344 4826 3372 6394
rect 3436 6322 3464 6598
rect 3507 6556 3815 6565
rect 3507 6554 3513 6556
rect 3569 6554 3593 6556
rect 3649 6554 3673 6556
rect 3729 6554 3753 6556
rect 3809 6554 3815 6556
rect 3569 6502 3571 6554
rect 3751 6502 3753 6554
rect 3507 6500 3513 6502
rect 3569 6500 3593 6502
rect 3649 6500 3673 6502
rect 3729 6500 3753 6502
rect 3809 6500 3815 6502
rect 3507 6491 3815 6500
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3507 5468 3815 5477
rect 3507 5466 3513 5468
rect 3569 5466 3593 5468
rect 3649 5466 3673 5468
rect 3729 5466 3753 5468
rect 3809 5466 3815 5468
rect 3569 5414 3571 5466
rect 3751 5414 3753 5466
rect 3507 5412 3513 5414
rect 3569 5412 3593 5414
rect 3649 5412 3673 5414
rect 3729 5412 3753 5414
rect 3809 5412 3815 5414
rect 3507 5403 3815 5412
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 2688 4694 2740 4700
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4214 2360 4422
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2056 3602 2084 4082
rect 2240 3738 2268 4150
rect 2700 4078 2728 4694
rect 3068 4678 3280 4706
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 3068 3942 3096 4678
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3252 4282 3280 4490
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3344 4214 3372 4762
rect 3507 4380 3815 4389
rect 3507 4378 3513 4380
rect 3569 4378 3593 4380
rect 3649 4378 3673 4380
rect 3729 4378 3753 4380
rect 3809 4378 3815 4380
rect 3569 4326 3571 4378
rect 3751 4326 3753 4378
rect 3507 4324 3513 4326
rect 3569 4324 3593 4326
rect 3649 4324 3673 4326
rect 3729 4324 3753 4326
rect 3809 4324 3815 4326
rect 3507 4315 3815 4324
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2847 3836 3155 3845
rect 2847 3834 2853 3836
rect 2909 3834 2933 3836
rect 2989 3834 3013 3836
rect 3069 3834 3093 3836
rect 3149 3834 3155 3836
rect 2909 3782 2911 3834
rect 3091 3782 3093 3834
rect 2847 3780 2853 3782
rect 2909 3780 2933 3782
rect 2989 3780 3013 3782
rect 3069 3780 3093 3782
rect 3149 3780 3155 3782
rect 2847 3771 3155 3780
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 3344 3534 3372 4150
rect 4172 4146 4200 4966
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4264 4078 4292 4558
rect 4356 4486 4384 9658
rect 4540 9654 4568 10066
rect 6380 9674 6408 11018
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 4528 9648 4580 9654
rect 6380 9646 6500 9674
rect 6564 9654 6592 10474
rect 6642 10364 6950 10373
rect 6642 10362 6648 10364
rect 6704 10362 6728 10364
rect 6784 10362 6808 10364
rect 6864 10362 6888 10364
rect 6944 10362 6950 10364
rect 6704 10310 6706 10362
rect 6886 10310 6888 10362
rect 6642 10308 6648 10310
rect 6704 10308 6728 10310
rect 6784 10308 6808 10310
rect 6864 10308 6888 10310
rect 6944 10308 6950 10310
rect 6642 10299 6950 10308
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 4528 9590 4580 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 8838 4568 9454
rect 5368 9178 5396 9522
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 9081 5488 9454
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5446 9072 5502 9081
rect 5828 9042 5856 9318
rect 5446 9007 5502 9016
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 6472 8906 6500 9646
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6932 9602 6960 9862
rect 7024 9704 7052 12038
rect 7208 11898 7236 12056
rect 7380 12038 7432 12044
rect 7302 11996 7610 12005
rect 7302 11994 7308 11996
rect 7364 11994 7388 11996
rect 7444 11994 7468 11996
rect 7524 11994 7548 11996
rect 7604 11994 7610 11996
rect 7364 11942 7366 11994
rect 7546 11942 7548 11994
rect 7302 11940 7308 11942
rect 7364 11940 7388 11942
rect 7444 11940 7468 11942
rect 7524 11940 7548 11942
rect 7604 11940 7610 11942
rect 7302 11931 7610 11940
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 10810 7236 11698
rect 7302 10908 7610 10917
rect 7302 10906 7308 10908
rect 7364 10906 7388 10908
rect 7444 10906 7468 10908
rect 7524 10906 7548 10908
rect 7604 10906 7610 10908
rect 7364 10854 7366 10906
rect 7546 10854 7548 10906
rect 7302 10852 7308 10854
rect 7364 10852 7388 10854
rect 7444 10852 7468 10854
rect 7524 10852 7548 10854
rect 7604 10852 7610 10854
rect 7302 10843 7610 10852
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7668 10674 7696 12406
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9926 7144 10406
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7208 9722 7236 10542
rect 7760 10266 7788 11290
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7302 9820 7610 9829
rect 7302 9818 7308 9820
rect 7364 9818 7388 9820
rect 7444 9818 7468 9820
rect 7524 9818 7548 9820
rect 7604 9818 7610 9820
rect 7364 9766 7366 9818
rect 7546 9766 7548 9818
rect 7302 9764 7308 9766
rect 7364 9764 7388 9766
rect 7444 9764 7468 9766
rect 7524 9764 7548 9766
rect 7604 9764 7610 9766
rect 7302 9755 7610 9764
rect 7668 9722 7696 9998
rect 7760 9926 7788 10066
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7104 9716 7156 9722
rect 7024 9676 7104 9704
rect 7104 9658 7156 9664
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 6932 9574 7052 9602
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9058 6592 9318
rect 6642 9276 6950 9285
rect 6642 9274 6648 9276
rect 6704 9274 6728 9276
rect 6784 9274 6808 9276
rect 6864 9274 6888 9276
rect 6944 9274 6950 9276
rect 6704 9222 6706 9274
rect 6886 9222 6888 9274
rect 6642 9220 6648 9222
rect 6704 9220 6728 9222
rect 6784 9220 6808 9222
rect 6864 9220 6888 9222
rect 6944 9220 6950 9222
rect 6642 9211 6950 9220
rect 6828 9104 6880 9110
rect 6564 9042 6776 9058
rect 6828 9046 6880 9052
rect 6564 9036 6788 9042
rect 6564 9030 6736 9036
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 7750 4568 8774
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7818 5304 8366
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4448 6662 4476 7278
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4436 6248 4488 6254
rect 4540 6236 4568 7686
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 4488 6208 4568 6236
rect 4712 6248 4764 6254
rect 4436 6190 4488 6196
rect 4712 6190 4764 6196
rect 4448 4826 4476 6190
rect 4724 5914 4752 6190
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5370 5856 5714
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5828 5114 5856 5170
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5736 5086 5856 5114
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 5184 4622 5212 5034
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4690 5672 4966
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3988 3534 4016 3878
rect 4264 3534 4292 4014
rect 4356 3738 4384 4082
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 3507 3292 3815 3301
rect 3507 3290 3513 3292
rect 3569 3290 3593 3292
rect 3649 3290 3673 3292
rect 3729 3290 3753 3292
rect 3809 3290 3815 3292
rect 3569 3238 3571 3290
rect 3751 3238 3753 3290
rect 3507 3236 3513 3238
rect 3569 3236 3593 3238
rect 3649 3236 3673 3238
rect 3729 3236 3753 3238
rect 3809 3236 3815 3238
rect 3507 3227 3815 3236
rect 4540 2774 4568 4558
rect 5276 3534 5304 4626
rect 5736 4486 5764 5086
rect 6012 4554 6040 7414
rect 6564 6866 6592 9030
rect 6736 8978 6788 8984
rect 6840 8634 6868 9046
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6642 8188 6950 8197
rect 6642 8186 6648 8188
rect 6704 8186 6728 8188
rect 6784 8186 6808 8188
rect 6864 8186 6888 8188
rect 6944 8186 6950 8188
rect 6704 8134 6706 8186
rect 6886 8134 6888 8186
rect 6642 8132 6648 8134
rect 6704 8132 6728 8134
rect 6784 8132 6808 8134
rect 6864 8132 6888 8134
rect 6944 8132 6950 8134
rect 6642 8123 6950 8132
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7546 6960 7686
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 7206 7052 9574
rect 7116 8566 7144 9658
rect 8036 9586 8064 12242
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11354 8248 12174
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11354 8432 12038
rect 8496 11830 8524 13874
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 12442 9904 13738
rect 9864 12436 9916 12442
rect 9784 12406 9864 12434
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10674 8248 10950
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8312 10266 8340 11154
rect 8496 11014 8524 11766
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11354 8616 11630
rect 9692 11558 9720 12174
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7208 8974 7236 9522
rect 8128 9382 8156 9862
rect 8220 9602 8248 9930
rect 8496 9926 8524 10134
rect 8772 9926 8800 10610
rect 9232 10266 9260 10678
rect 9220 10260 9272 10266
rect 9140 10220 9220 10248
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9704 8800 9862
rect 8588 9676 8800 9704
rect 8300 9648 8352 9654
rect 8220 9596 8300 9602
rect 8220 9590 8352 9596
rect 8220 9574 8340 9590
rect 8588 9586 8616 9676
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9058 8156 9318
rect 8036 9030 8156 9058
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7302 8732 7610 8741
rect 7302 8730 7308 8732
rect 7364 8730 7388 8732
rect 7444 8730 7468 8732
rect 7524 8730 7548 8732
rect 7604 8730 7610 8732
rect 7364 8678 7366 8730
rect 7546 8678 7548 8730
rect 7302 8676 7308 8678
rect 7364 8676 7388 8678
rect 7444 8676 7468 8678
rect 7524 8676 7548 8678
rect 7604 8676 7610 8678
rect 7302 8667 7610 8676
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7760 8362 7788 8842
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7302 7644 7610 7653
rect 7302 7642 7308 7644
rect 7364 7642 7388 7644
rect 7444 7642 7468 7644
rect 7524 7642 7548 7644
rect 7604 7642 7610 7644
rect 7364 7590 7366 7642
rect 7546 7590 7548 7642
rect 7302 7588 7308 7590
rect 7364 7588 7388 7590
rect 7444 7588 7468 7590
rect 7524 7588 7548 7590
rect 7604 7588 7610 7590
rect 7302 7579 7610 7588
rect 7760 7546 7788 8298
rect 8036 8090 8064 9030
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8634 8156 8910
rect 8220 8634 8248 9454
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8378 8340 9574
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8404 9178 8432 9522
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8496 8498 8524 9386
rect 8588 9042 8616 9522
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8680 8974 8708 9522
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8220 8350 8340 8378
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8220 7886 8248 8350
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8404 7546 8432 8230
rect 8496 8090 8524 8434
rect 9140 8090 9168 10220
rect 9220 10202 9272 10208
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9178 9260 9998
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 8362 9260 8774
rect 9324 8634 9352 11086
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9416 10044 9444 10610
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9692 10130 9720 11494
rect 9784 11218 9812 12406
rect 9864 12378 9916 12384
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9784 10742 9812 11018
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9496 10056 9548 10062
rect 9416 10016 9496 10044
rect 9496 9998 9548 10004
rect 9508 9586 9536 9998
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 8922 9536 9522
rect 9784 9178 9812 10066
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9586 9072 9642 9081
rect 9586 9007 9588 9016
rect 9640 9007 9642 9016
rect 9680 9036 9732 9042
rect 9588 8978 9640 8984
rect 9680 8978 9732 8984
rect 9692 8922 9720 8978
rect 9508 8894 9720 8922
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9232 7750 9260 8298
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6642 7100 6950 7109
rect 6642 7098 6648 7100
rect 6704 7098 6728 7100
rect 6784 7098 6808 7100
rect 6864 7098 6888 7100
rect 6944 7098 6950 7100
rect 6704 7046 6706 7098
rect 6886 7046 6888 7098
rect 6642 7044 6648 7046
rect 6704 7044 6728 7046
rect 6784 7044 6808 7046
rect 6864 7044 6888 7046
rect 6944 7044 6950 7046
rect 6642 7035 6950 7044
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 5778 6316 6734
rect 7208 6730 7236 7278
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6254 6500 6598
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5914 6408 6054
rect 6642 6012 6950 6021
rect 6642 6010 6648 6012
rect 6704 6010 6728 6012
rect 6784 6010 6808 6012
rect 6864 6010 6888 6012
rect 6944 6010 6950 6012
rect 6704 5958 6706 6010
rect 6886 5958 6888 6010
rect 6642 5956 6648 5958
rect 6704 5956 6728 5958
rect 6784 5956 6808 5958
rect 6864 5956 6888 5958
rect 6944 5956 6950 5958
rect 6642 5947 6950 5956
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 7208 5846 7236 6666
rect 7302 6556 7610 6565
rect 7302 6554 7308 6556
rect 7364 6554 7388 6556
rect 7444 6554 7468 6556
rect 7524 6554 7548 6556
rect 7604 6554 7610 6556
rect 7364 6502 7366 6554
rect 7546 6502 7548 6554
rect 7302 6500 7308 6502
rect 7364 6500 7388 6502
rect 7444 6500 7468 6502
rect 7524 6500 7548 6502
rect 7604 6500 7610 6502
rect 7302 6491 7610 6500
rect 8956 6458 8984 7278
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9232 6390 9260 7686
rect 9416 7546 9444 8230
rect 9876 8090 9904 11766
rect 9968 11762 9996 14282
rect 10060 13802 10088 14436
rect 10232 14418 10284 14424
rect 10336 13938 10364 14486
rect 10796 14074 10824 15302
rect 10980 15042 11008 15302
rect 11097 15260 11405 15269
rect 11097 15258 11103 15260
rect 11159 15258 11183 15260
rect 11239 15258 11263 15260
rect 11319 15258 11343 15260
rect 11399 15258 11405 15260
rect 11159 15206 11161 15258
rect 11341 15206 11343 15258
rect 11097 15204 11103 15206
rect 11159 15204 11183 15206
rect 11239 15204 11263 15206
rect 11319 15204 11343 15206
rect 11399 15204 11405 15206
rect 11097 15195 11405 15204
rect 10980 15014 11100 15042
rect 11072 14414 11100 15014
rect 11440 14890 11468 15302
rect 11532 14958 11560 15438
rect 11624 15162 11652 15982
rect 14232 15804 14540 15813
rect 14232 15802 14238 15804
rect 14294 15802 14318 15804
rect 14374 15802 14398 15804
rect 14454 15802 14478 15804
rect 14534 15802 14540 15804
rect 14294 15750 14296 15802
rect 14476 15750 14478 15802
rect 14232 15748 14238 15750
rect 14294 15748 14318 15750
rect 14374 15748 14398 15750
rect 14454 15748 14478 15750
rect 14534 15748 14540 15750
rect 14232 15739 14540 15748
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11808 15450 11836 15574
rect 14648 15496 14700 15502
rect 11808 15422 11928 15450
rect 14648 15438 14700 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11532 14414 11560 14894
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11097 14172 11405 14181
rect 11097 14170 11103 14172
rect 11159 14170 11183 14172
rect 11239 14170 11263 14172
rect 11319 14170 11343 14172
rect 11399 14170 11405 14172
rect 11159 14118 11161 14170
rect 11341 14118 11343 14170
rect 11097 14116 11103 14118
rect 11159 14116 11183 14118
rect 11239 14116 11263 14118
rect 11319 14116 11343 14118
rect 11399 14116 11405 14118
rect 11097 14107 11405 14116
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10437 13628 10745 13637
rect 10437 13626 10443 13628
rect 10499 13626 10523 13628
rect 10579 13626 10603 13628
rect 10659 13626 10683 13628
rect 10739 13626 10745 13628
rect 10499 13574 10501 13626
rect 10681 13574 10683 13626
rect 10437 13572 10443 13574
rect 10499 13572 10523 13574
rect 10579 13572 10603 13574
rect 10659 13572 10683 13574
rect 10739 13572 10745 13574
rect 10437 13563 10745 13572
rect 11097 13084 11405 13093
rect 11097 13082 11103 13084
rect 11159 13082 11183 13084
rect 11239 13082 11263 13084
rect 11319 13082 11343 13084
rect 11399 13082 11405 13084
rect 11159 13030 11161 13082
rect 11341 13030 11343 13082
rect 11097 13028 11103 13030
rect 11159 13028 11183 13030
rect 11239 13028 11263 13030
rect 11319 13028 11343 13030
rect 11399 13028 11405 13030
rect 11097 13019 11405 13028
rect 11532 12850 11560 14350
rect 11808 14074 11836 15302
rect 11900 14414 11928 15422
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14074 11928 14214
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 12084 13530 12112 15370
rect 12544 15162 12572 15370
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12544 14414 12572 15098
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 14074 12204 14214
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 11900 12986 11928 13126
rect 12452 12986 12480 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12918 12572 14350
rect 12820 14006 12848 14758
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12808 14000 12860 14006
rect 13096 13954 13124 14962
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12808 13942 12860 13948
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12728 13818 12756 13942
rect 13004 13926 13124 13954
rect 13004 13870 13032 13926
rect 12992 13864 13044 13870
rect 12636 13394 12664 13806
rect 12728 13802 12848 13818
rect 12992 13806 13044 13812
rect 12728 13796 12860 13802
rect 12728 13790 12808 13796
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 10437 12540 10745 12549
rect 10437 12538 10443 12540
rect 10499 12538 10523 12540
rect 10579 12538 10603 12540
rect 10659 12538 10683 12540
rect 10739 12538 10745 12540
rect 10499 12486 10501 12538
rect 10681 12486 10683 12538
rect 10437 12484 10443 12486
rect 10499 12484 10523 12486
rect 10579 12484 10603 12486
rect 10659 12484 10683 12486
rect 10739 12484 10745 12486
rect 10437 12475 10745 12484
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11898 10732 12038
rect 11097 11996 11405 12005
rect 11097 11994 11103 11996
rect 11159 11994 11183 11996
rect 11239 11994 11263 11996
rect 11319 11994 11343 11996
rect 11399 11994 11405 11996
rect 11159 11942 11161 11994
rect 11341 11942 11343 11994
rect 11097 11940 11103 11942
rect 11159 11940 11183 11942
rect 11239 11940 11263 11942
rect 11319 11940 11343 11942
rect 11399 11940 11405 11942
rect 11097 11931 11405 11940
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 11532 11694 11560 12786
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 9926 9996 10950
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 10060 8974 10088 10406
rect 10152 10266 10180 11086
rect 10336 10742 10364 11494
rect 10437 11452 10745 11461
rect 10437 11450 10443 11452
rect 10499 11450 10523 11452
rect 10579 11450 10603 11452
rect 10659 11450 10683 11452
rect 10739 11450 10745 11452
rect 10499 11398 10501 11450
rect 10681 11398 10683 11450
rect 10437 11396 10443 11398
rect 10499 11396 10523 11398
rect 10579 11396 10603 11398
rect 10659 11396 10683 11398
rect 10739 11396 10745 11398
rect 10437 11387 10745 11396
rect 10888 11354 10916 11494
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10437 10364 10745 10373
rect 10437 10362 10443 10364
rect 10499 10362 10523 10364
rect 10579 10362 10603 10364
rect 10659 10362 10683 10364
rect 10739 10362 10745 10364
rect 10499 10310 10501 10362
rect 10681 10310 10683 10362
rect 10437 10308 10443 10310
rect 10499 10308 10523 10310
rect 10579 10308 10603 10310
rect 10659 10308 10683 10310
rect 10739 10308 10745 10310
rect 10437 10299 10745 10308
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10980 10062 11008 11290
rect 11532 11218 11560 11630
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11808 11150 11836 12038
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11097 10908 11405 10917
rect 11097 10906 11103 10908
rect 11159 10906 11183 10908
rect 11239 10906 11263 10908
rect 11319 10906 11343 10908
rect 11399 10906 11405 10908
rect 11159 10854 11161 10906
rect 11341 10854 11343 10906
rect 11097 10852 11103 10854
rect 11159 10852 11183 10854
rect 11239 10852 11263 10854
rect 11319 10852 11343 10854
rect 11399 10852 11405 10854
rect 11097 10843 11405 10852
rect 11440 10742 11468 10950
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10336 9722 10364 9998
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10612 9722 10640 9930
rect 11097 9820 11405 9829
rect 11097 9818 11103 9820
rect 11159 9818 11183 9820
rect 11239 9818 11263 9820
rect 11319 9818 11343 9820
rect 11399 9818 11405 9820
rect 11159 9766 11161 9818
rect 11341 9766 11343 9818
rect 11097 9764 11103 9766
rect 11159 9764 11183 9766
rect 11239 9764 11263 9766
rect 11319 9764 11343 9766
rect 11399 9764 11405 9766
rect 11097 9755 11405 9764
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10152 8498 10180 9454
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8634 10272 8910
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9508 7562 9536 8026
rect 9876 7834 9904 8026
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9784 7806 9904 7834
rect 9600 7698 9628 7754
rect 9600 7670 9720 7698
rect 9404 7540 9456 7546
rect 9508 7534 9628 7562
rect 9404 7482 9456 7488
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6748 5166 6776 5714
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 5012 6776 5102
rect 6564 4984 6776 5012
rect 6564 4826 6592 4984
rect 6642 4924 6950 4933
rect 6642 4922 6648 4924
rect 6704 4922 6728 4924
rect 6784 4922 6808 4924
rect 6864 4922 6888 4924
rect 6944 4922 6950 4924
rect 6704 4870 6706 4922
rect 6886 4870 6888 4922
rect 6642 4868 6648 4870
rect 6704 4868 6728 4870
rect 6784 4868 6808 4870
rect 6864 4868 6888 4870
rect 6944 4868 6950 4870
rect 6642 4859 6950 4868
rect 7208 4826 7236 5646
rect 7302 5468 7610 5477
rect 7302 5466 7308 5468
rect 7364 5466 7388 5468
rect 7444 5466 7468 5468
rect 7524 5466 7548 5468
rect 7604 5466 7610 5468
rect 7364 5414 7366 5466
rect 7546 5414 7548 5466
rect 7302 5412 7308 5414
rect 7364 5412 7388 5414
rect 7444 5412 7468 5414
rect 7524 5412 7548 5414
rect 7604 5412 7610 5414
rect 7302 5403 7610 5412
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4826 8708 4966
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4146 5764 4422
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5920 3942 5948 4082
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5736 3058 5764 3402
rect 5828 3194 5856 3878
rect 5920 3738 5948 3878
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6012 3466 6040 4490
rect 7208 4146 7236 4762
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7302 4380 7610 4389
rect 7302 4378 7308 4380
rect 7364 4378 7388 4380
rect 7444 4378 7468 4380
rect 7524 4378 7548 4380
rect 7604 4378 7610 4380
rect 7364 4326 7366 4378
rect 7546 4326 7548 4378
rect 7302 4324 7308 4326
rect 7364 4324 7388 4326
rect 7444 4324 7468 4326
rect 7524 4324 7548 4326
rect 7604 4324 7610 4326
rect 7302 4315 7610 4324
rect 8128 4146 8156 4422
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6104 3738 6132 4014
rect 6642 3836 6950 3845
rect 6642 3834 6648 3836
rect 6704 3834 6728 3836
rect 6784 3834 6808 3836
rect 6864 3834 6888 3836
rect 6944 3834 6950 3836
rect 6704 3782 6706 3834
rect 6886 3782 6888 3834
rect 6642 3780 6648 3782
rect 6704 3780 6728 3782
rect 6784 3780 6808 3782
rect 6864 3780 6888 3782
rect 6944 3780 6950 3782
rect 6642 3771 6950 3780
rect 7208 3738 7236 4082
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 8128 3534 8156 4082
rect 8220 3534 8248 4490
rect 9048 4282 9076 5306
rect 9416 5234 9444 7142
rect 9600 6066 9628 7534
rect 9692 6254 9720 7670
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 6186 9812 7806
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 6866 9904 7686
rect 9968 7546 9996 8366
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9600 6038 9812 6066
rect 9784 5710 9812 6038
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9763 5704 9815 5710
rect 9763 5646 9815 5652
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9140 4282 9168 4626
rect 9232 4486 9260 4966
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8680 3738 8708 3878
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 9140 3602 9168 4218
rect 9508 4078 9536 5646
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5370 9628 5510
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9678 5264 9734 5273
rect 9588 5228 9640 5234
rect 9678 5199 9680 5208
rect 9588 5170 9640 5176
rect 9732 5199 9734 5208
rect 9680 5170 9732 5176
rect 9600 4486 9628 5170
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9600 4026 9628 4422
rect 9692 4146 9720 4966
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9600 3998 9720 4026
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6748 3126 6776 3334
rect 7302 3292 7610 3301
rect 7302 3290 7308 3292
rect 7364 3290 7388 3292
rect 7444 3290 7468 3292
rect 7524 3290 7548 3292
rect 7604 3290 7610 3292
rect 7364 3238 7366 3290
rect 7546 3238 7548 3290
rect 7302 3236 7308 3238
rect 7364 3236 7388 3238
rect 7444 3236 7468 3238
rect 7524 3236 7548 3238
rect 7604 3236 7610 3238
rect 7302 3227 7610 3236
rect 8128 3194 8156 3470
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 8220 3058 8248 3470
rect 9600 3466 9628 3538
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9692 3194 9720 3998
rect 9784 3942 9812 5646
rect 9876 4554 9904 6258
rect 9968 5302 9996 6258
rect 10152 5914 10180 6326
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 5370 10088 5646
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10152 5216 10180 5850
rect 10336 5710 10364 9658
rect 10506 9616 10562 9625
rect 11808 9586 11836 11086
rect 12360 10674 12388 11630
rect 12544 11150 12572 12854
rect 12636 12306 12664 13330
rect 12728 13258 12756 13790
rect 12808 13738 12860 13744
rect 13372 13530 13400 14758
rect 13832 14618 13860 15030
rect 14016 15026 14044 15302
rect 14108 15162 14136 15302
rect 14660 15162 14688 15438
rect 14892 15260 15200 15269
rect 14892 15258 14898 15260
rect 14954 15258 14978 15260
rect 15034 15258 15058 15260
rect 15114 15258 15138 15260
rect 15194 15258 15200 15260
rect 14954 15206 14956 15258
rect 15136 15206 15138 15258
rect 14892 15204 14898 15206
rect 14954 15204 14978 15206
rect 15034 15204 15058 15206
rect 15114 15204 15138 15206
rect 15194 15204 15200 15206
rect 14892 15195 15200 15204
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14232 14716 14540 14725
rect 14232 14714 14238 14716
rect 14294 14714 14318 14716
rect 14374 14714 14398 14716
rect 14454 14714 14478 14716
rect 14534 14714 14540 14716
rect 14294 14662 14296 14714
rect 14476 14662 14478 14714
rect 14232 14660 14238 14662
rect 14294 14660 14318 14662
rect 14374 14660 14398 14662
rect 14454 14660 14478 14662
rect 14534 14660 14540 14662
rect 14232 14651 14540 14660
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 14074 13676 14282
rect 14892 14172 15200 14181
rect 14892 14170 14898 14172
rect 14954 14170 14978 14172
rect 15034 14170 15058 14172
rect 15114 14170 15138 14172
rect 15194 14170 15200 14172
rect 14954 14118 14956 14170
rect 15136 14118 15138 14170
rect 14892 14116 14898 14118
rect 14954 14116 14978 14118
rect 15034 14116 15058 14118
rect 15114 14116 15138 14118
rect 15194 14116 15200 14118
rect 14892 14107 15200 14116
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 14232 13628 14540 13637
rect 14232 13626 14238 13628
rect 14294 13626 14318 13628
rect 14374 13626 14398 13628
rect 14454 13626 14478 13628
rect 14534 13626 14540 13628
rect 14294 13574 14296 13626
rect 14476 13574 14478 13626
rect 14232 13572 14238 13574
rect 14294 13572 14318 13574
rect 14374 13572 14398 13574
rect 14454 13572 14478 13574
rect 14534 13572 14540 13574
rect 14232 13563 14540 13572
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 14892 13084 15200 13093
rect 14892 13082 14898 13084
rect 14954 13082 14978 13084
rect 15034 13082 15058 13084
rect 15114 13082 15138 13084
rect 15194 13082 15200 13084
rect 14954 13030 14956 13082
rect 15136 13030 15138 13082
rect 14892 13028 14898 13030
rect 14954 13028 14978 13030
rect 15034 13028 15058 13030
rect 15114 13028 15138 13030
rect 15194 13028 15200 13030
rect 14892 13019 15200 13028
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 13372 12238 13400 12582
rect 14232 12540 14540 12549
rect 14232 12538 14238 12540
rect 14294 12538 14318 12540
rect 14374 12538 14398 12540
rect 14454 12538 14478 12540
rect 14534 12538 14540 12540
rect 14294 12486 14296 12538
rect 14476 12486 14478 12538
rect 14232 12484 14238 12486
rect 14294 12484 14318 12486
rect 14374 12484 14398 12486
rect 14454 12484 14478 12486
rect 14534 12484 14540 12486
rect 14232 12475 14540 12484
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12636 11354 12664 11698
rect 13556 11694 13584 12038
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 13556 11218 13584 11630
rect 14232 11452 14540 11461
rect 14232 11450 14238 11452
rect 14294 11450 14318 11452
rect 14374 11450 14398 11452
rect 14454 11450 14478 11452
rect 14534 11450 14540 11452
rect 14294 11398 14296 11450
rect 14476 11398 14478 11450
rect 14232 11396 14238 11398
rect 14294 11396 14318 11398
rect 14374 11396 14398 11398
rect 14454 11396 14478 11398
rect 14534 11396 14540 11398
rect 14232 11387 14540 11396
rect 14568 11354 14596 12038
rect 14660 11898 14688 12174
rect 14752 11898 14780 12174
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14892 11996 15200 12005
rect 14892 11994 14898 11996
rect 14954 11994 14978 11996
rect 15034 11994 15058 11996
rect 15114 11994 15138 11996
rect 15194 11994 15200 11996
rect 14954 11942 14956 11994
rect 15136 11942 15138 11994
rect 14892 11940 14898 11942
rect 14954 11940 14978 11942
rect 15034 11940 15058 11942
rect 15114 11940 15138 11942
rect 15194 11940 15200 11942
rect 14892 11931 15200 11940
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 15304 11830 15332 12038
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10742 13768 11086
rect 13832 10742 13860 11222
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 12360 10266 12388 10610
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 10506 9551 10508 9560
rect 10560 9551 10562 9560
rect 10876 9580 10928 9586
rect 10508 9522 10560 9528
rect 10876 9522 10928 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 10437 9276 10745 9285
rect 10437 9274 10443 9276
rect 10499 9274 10523 9276
rect 10579 9274 10603 9276
rect 10659 9274 10683 9276
rect 10739 9274 10745 9276
rect 10499 9222 10501 9274
rect 10681 9222 10683 9274
rect 10437 9220 10443 9222
rect 10499 9220 10523 9222
rect 10579 9220 10603 9222
rect 10659 9220 10683 9222
rect 10739 9220 10745 9222
rect 10437 9211 10745 9220
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8566 10640 8774
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10704 8514 10732 8910
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10796 8634 10824 8842
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10704 8486 10824 8514
rect 10437 8188 10745 8197
rect 10437 8186 10443 8188
rect 10499 8186 10523 8188
rect 10579 8186 10603 8188
rect 10659 8186 10683 8188
rect 10739 8186 10745 8188
rect 10499 8134 10501 8186
rect 10681 8134 10683 8186
rect 10437 8132 10443 8134
rect 10499 8132 10523 8134
rect 10579 8132 10603 8134
rect 10659 8132 10683 8134
rect 10739 8132 10745 8134
rect 10437 8123 10745 8132
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10704 7750 10732 8026
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10437 7100 10745 7109
rect 10437 7098 10443 7100
rect 10499 7098 10523 7100
rect 10579 7098 10603 7100
rect 10659 7098 10683 7100
rect 10739 7098 10745 7100
rect 10499 7046 10501 7098
rect 10681 7046 10683 7098
rect 10437 7044 10443 7046
rect 10499 7044 10523 7046
rect 10579 7044 10603 7046
rect 10659 7044 10683 7046
rect 10739 7044 10745 7046
rect 10437 7035 10745 7044
rect 10437 6012 10745 6021
rect 10437 6010 10443 6012
rect 10499 6010 10523 6012
rect 10579 6010 10603 6012
rect 10659 6010 10683 6012
rect 10739 6010 10745 6012
rect 10499 5958 10501 6010
rect 10681 5958 10683 6010
rect 10437 5956 10443 5958
rect 10499 5956 10523 5958
rect 10579 5956 10603 5958
rect 10659 5956 10683 5958
rect 10739 5956 10745 5958
rect 10437 5947 10745 5956
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10060 5188 10180 5216
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 4282 9904 4490
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9876 3398 9904 4218
rect 10060 3602 10088 5188
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 3738 10180 5034
rect 10428 5030 10456 5102
rect 10796 5030 10824 8486
rect 10888 8090 10916 9522
rect 13464 9518 13492 10610
rect 13924 10266 13952 11018
rect 14232 10364 14540 10373
rect 14232 10362 14238 10364
rect 14294 10362 14318 10364
rect 14374 10362 14398 10364
rect 14454 10362 14478 10364
rect 14534 10362 14540 10364
rect 14294 10310 14296 10362
rect 14476 10310 14478 10362
rect 14232 10308 14238 10310
rect 14294 10308 14318 10310
rect 14374 10308 14398 10310
rect 14454 10308 14478 10310
rect 14534 10308 14540 10310
rect 14232 10299 14540 10308
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14108 9722 14136 10134
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10980 8634 11008 9318
rect 11256 8906 11284 9318
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 11097 8732 11405 8741
rect 11097 8730 11103 8732
rect 11159 8730 11183 8732
rect 11239 8730 11263 8732
rect 11319 8730 11343 8732
rect 11399 8730 11405 8732
rect 11159 8678 11161 8730
rect 11341 8678 11343 8730
rect 11097 8676 11103 8678
rect 11159 8676 11183 8678
rect 11239 8676 11263 8678
rect 11319 8676 11343 8678
rect 11399 8676 11405 8678
rect 11097 8667 11405 8676
rect 12912 8634 12940 8774
rect 13464 8634 13492 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10888 6866 10916 8026
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10980 6458 11008 8230
rect 11097 7644 11405 7653
rect 11097 7642 11103 7644
rect 11159 7642 11183 7644
rect 11239 7642 11263 7644
rect 11319 7642 11343 7644
rect 11399 7642 11405 7644
rect 11159 7590 11161 7642
rect 11341 7590 11343 7642
rect 11097 7588 11103 7590
rect 11159 7588 11183 7590
rect 11239 7588 11263 7590
rect 11319 7588 11343 7590
rect 11399 7588 11405 7590
rect 11097 7579 11405 7588
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6798 11192 7142
rect 11256 7002 11284 7414
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11097 6556 11405 6565
rect 11097 6554 11103 6556
rect 11159 6554 11183 6556
rect 11239 6554 11263 6556
rect 11319 6554 11343 6556
rect 11399 6554 11405 6556
rect 11159 6502 11161 6554
rect 11341 6502 11343 6554
rect 11097 6500 11103 6502
rect 11159 6500 11183 6502
rect 11239 6500 11263 6502
rect 11319 6500 11343 6502
rect 11399 6500 11405 6502
rect 11097 6491 11405 6500
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10437 4924 10745 4933
rect 10437 4922 10443 4924
rect 10499 4922 10523 4924
rect 10579 4922 10603 4924
rect 10659 4922 10683 4924
rect 10739 4922 10745 4924
rect 10499 4870 10501 4922
rect 10681 4870 10683 4922
rect 10437 4868 10443 4870
rect 10499 4868 10523 4870
rect 10579 4868 10603 4870
rect 10659 4868 10683 4870
rect 10739 4868 10745 4870
rect 10437 4859 10745 4868
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4282 10824 4490
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10437 3836 10745 3845
rect 10437 3834 10443 3836
rect 10499 3834 10523 3836
rect 10579 3834 10603 3836
rect 10659 3834 10683 3836
rect 10739 3834 10745 3836
rect 10499 3782 10501 3834
rect 10681 3782 10683 3834
rect 10437 3780 10443 3782
rect 10499 3780 10523 3782
rect 10579 3780 10603 3782
rect 10659 3780 10683 3782
rect 10739 3780 10745 3782
rect 10437 3771 10745 3780
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3194 9904 3334
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10888 3058 10916 6054
rect 10980 5710 11008 6394
rect 11440 6390 11468 8502
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7818 11560 8230
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11716 6662 11744 8434
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7954 12296 8230
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 7410 12020 7822
rect 12820 7546 12848 8366
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13280 8090 13308 8298
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13832 7750 13860 9454
rect 14232 9276 14540 9285
rect 14232 9274 14238 9276
rect 14294 9274 14318 9276
rect 14374 9274 14398 9276
rect 14454 9274 14478 9276
rect 14534 9274 14540 9276
rect 14294 9222 14296 9274
rect 14476 9222 14478 9274
rect 14232 9220 14238 9222
rect 14294 9220 14318 9222
rect 14374 9220 14398 9222
rect 14454 9220 14478 9222
rect 14534 9220 14540 9222
rect 14232 9211 14540 9220
rect 14568 9178 14596 10066
rect 14660 10062 14688 11494
rect 14752 11014 14780 11698
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11218 15424 11630
rect 15856 11354 15884 12174
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10690 14780 10950
rect 14892 10908 15200 10917
rect 14892 10906 14898 10908
rect 14954 10906 14978 10908
rect 15034 10906 15058 10908
rect 15114 10906 15138 10908
rect 15194 10906 15200 10908
rect 14954 10854 14956 10906
rect 15136 10854 15138 10906
rect 14892 10852 14898 10854
rect 14954 10852 14978 10854
rect 15034 10852 15058 10854
rect 15114 10852 15138 10854
rect 15194 10852 15200 10854
rect 14892 10843 15200 10852
rect 14752 10674 14872 10690
rect 14752 10668 14884 10674
rect 14752 10662 14832 10668
rect 14832 10610 14884 10616
rect 14648 10056 14700 10062
rect 14844 10010 14872 10610
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14648 9998 14700 10004
rect 14752 9982 14872 10010
rect 14752 9518 14780 9982
rect 14892 9820 15200 9829
rect 14892 9818 14898 9820
rect 14954 9818 14978 9820
rect 15034 9818 15058 9820
rect 15114 9818 15138 9820
rect 15194 9818 15200 9820
rect 14954 9766 14956 9818
rect 15136 9766 15138 9818
rect 14892 9764 14898 9766
rect 14954 9764 14978 9766
rect 15034 9764 15058 9766
rect 15114 9764 15138 9766
rect 15194 9764 15200 9766
rect 14892 9755 15200 9764
rect 15304 9586 15332 10406
rect 15396 10266 15424 11154
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15488 9722 15516 9862
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14016 7546 14044 8502
rect 14200 8430 14228 8978
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14292 8634 14320 8842
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14108 8090 14136 8230
rect 14232 8188 14540 8197
rect 14232 8186 14238 8188
rect 14294 8186 14318 8188
rect 14374 8186 14398 8188
rect 14454 8186 14478 8188
rect 14534 8186 14540 8188
rect 14294 8134 14296 8186
rect 14476 8134 14478 8186
rect 14232 8132 14238 8134
rect 14294 8132 14318 8134
rect 14374 8132 14398 8134
rect 14454 8132 14478 8134
rect 14534 8132 14540 8134
rect 14232 8123 14540 8132
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 6866 12020 7346
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11992 5914 12020 6802
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10980 5166 11008 5646
rect 11097 5468 11405 5477
rect 11097 5466 11103 5468
rect 11159 5466 11183 5468
rect 11239 5466 11263 5468
rect 11319 5466 11343 5468
rect 11399 5466 11405 5468
rect 11159 5414 11161 5466
rect 11341 5414 11343 5466
rect 11097 5412 11103 5414
rect 11159 5412 11183 5414
rect 11239 5412 11263 5414
rect 11319 5412 11343 5414
rect 11399 5412 11405 5414
rect 11097 5403 11405 5412
rect 11336 5296 11388 5302
rect 11334 5264 11336 5273
rect 11388 5264 11390 5273
rect 11334 5199 11390 5208
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 10980 4826 11008 5102
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11348 4486 11376 5102
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4826 11468 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11992 4690 12020 5850
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12084 5234 12112 5510
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11097 4380 11405 4389
rect 11097 4378 11103 4380
rect 11159 4378 11183 4380
rect 11239 4378 11263 4380
rect 11319 4378 11343 4380
rect 11399 4378 11405 4380
rect 11159 4326 11161 4378
rect 11341 4326 11343 4378
rect 11097 4324 11103 4326
rect 11159 4324 11183 4326
rect 11239 4324 11263 4326
rect 11319 4324 11343 4326
rect 11399 4324 11405 4326
rect 11097 4315 11405 4324
rect 11992 4146 12020 4626
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11072 3738 11100 4014
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 3194 11008 3538
rect 11097 3292 11405 3301
rect 11097 3290 11103 3292
rect 11159 3290 11183 3292
rect 11239 3290 11263 3292
rect 11319 3290 11343 3292
rect 11399 3290 11405 3292
rect 11159 3238 11161 3290
rect 11341 3238 11343 3290
rect 11097 3236 11103 3238
rect 11159 3236 11183 3238
rect 11239 3236 11263 3238
rect 11319 3236 11343 3238
rect 11399 3236 11405 3238
rect 11097 3227 11405 3236
rect 11440 3194 11468 3946
rect 12636 3942 12664 5170
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3738 12664 3878
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 12636 3058 12664 3674
rect 12728 3534 12756 4422
rect 12820 4078 12848 4966
rect 12912 4622 12940 7482
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13924 7002 13952 7278
rect 14108 7206 14136 7822
rect 14660 7342 14688 8230
rect 14752 7546 14780 8774
rect 14892 8732 15200 8741
rect 14892 8730 14898 8732
rect 14954 8730 14978 8732
rect 15034 8730 15058 8732
rect 15114 8730 15138 8732
rect 15194 8730 15200 8732
rect 14954 8678 14956 8730
rect 15136 8678 15138 8730
rect 14892 8676 14898 8678
rect 14954 8676 14978 8678
rect 15034 8676 15058 8678
rect 15114 8676 15138 8678
rect 15194 8676 15200 8678
rect 14892 8667 15200 8676
rect 15304 8634 15332 9318
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 14892 7644 15200 7653
rect 14892 7642 14898 7644
rect 14954 7642 14978 7644
rect 15034 7642 15058 7644
rect 15114 7642 15138 7644
rect 15194 7642 15200 7644
rect 14954 7590 14956 7642
rect 15136 7590 15138 7642
rect 14892 7588 14898 7590
rect 14954 7588 14978 7590
rect 15034 7588 15058 7590
rect 15114 7588 15138 7590
rect 15194 7588 15200 7590
rect 14892 7579 15200 7588
rect 15396 7546 15424 9046
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 8294 15516 8910
rect 15580 8634 15608 9862
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 14108 6866 14136 7142
rect 14232 7100 14540 7109
rect 14232 7098 14238 7100
rect 14294 7098 14318 7100
rect 14374 7098 14398 7100
rect 14454 7098 14478 7100
rect 14534 7098 14540 7100
rect 14294 7046 14296 7098
rect 14476 7046 14478 7098
rect 14232 7044 14238 7046
rect 14294 7044 14318 7046
rect 14374 7044 14398 7046
rect 14454 7044 14478 7046
rect 14534 7044 14540 7046
rect 14232 7035 14540 7044
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14660 6730 14688 7142
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14232 6012 14540 6021
rect 14232 6010 14238 6012
rect 14294 6010 14318 6012
rect 14374 6010 14398 6012
rect 14454 6010 14478 6012
rect 14534 6010 14540 6012
rect 14294 5958 14296 6010
rect 14476 5958 14478 6010
rect 14232 5956 14238 5958
rect 14294 5956 14318 5958
rect 14374 5956 14398 5958
rect 14454 5956 14478 5958
rect 14534 5956 14540 5958
rect 14232 5947 14540 5956
rect 14752 5914 14780 7482
rect 15384 7336 15436 7342
rect 15488 7290 15516 7822
rect 15436 7284 15516 7290
rect 15384 7278 15516 7284
rect 15396 7262 15516 7278
rect 15396 6798 15424 7262
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15488 7002 15516 7142
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 14892 6556 15200 6565
rect 14892 6554 14898 6556
rect 14954 6554 14978 6556
rect 15034 6554 15058 6556
rect 15114 6554 15138 6556
rect 15194 6554 15200 6556
rect 14954 6502 14956 6554
rect 15136 6502 15138 6554
rect 14892 6500 14898 6502
rect 14954 6500 14978 6502
rect 15034 6500 15058 6502
rect 15114 6500 15138 6502
rect 15194 6500 15200 6502
rect 14892 6491 15200 6500
rect 15672 6458 15700 8978
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15856 8090 15884 8298
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15856 7426 15884 8026
rect 15764 7398 15884 7426
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6322 15792 7398
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15856 5914 15884 6598
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 14892 5468 15200 5477
rect 14892 5466 14898 5468
rect 14954 5466 14978 5468
rect 15034 5466 15058 5468
rect 15114 5466 15138 5468
rect 15194 5466 15200 5468
rect 14954 5414 14956 5466
rect 15136 5414 15138 5466
rect 14892 5412 14898 5414
rect 14954 5412 14978 5414
rect 15034 5412 15058 5414
rect 15114 5412 15138 5414
rect 15194 5412 15200 5414
rect 14892 5403 15200 5412
rect 14232 4924 14540 4933
rect 14232 4922 14238 4924
rect 14294 4922 14318 4924
rect 14374 4922 14398 4924
rect 14454 4922 14478 4924
rect 14534 4922 14540 4924
rect 14294 4870 14296 4922
rect 14476 4870 14478 4922
rect 14232 4868 14238 4870
rect 14294 4868 14318 4870
rect 14374 4868 14398 4870
rect 14454 4868 14478 4870
rect 14534 4868 14540 4870
rect 14232 4859 14540 4868
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12912 4214 12940 4558
rect 14892 4380 15200 4389
rect 14892 4378 14898 4380
rect 14954 4378 14978 4380
rect 15034 4378 15058 4380
rect 15114 4378 15138 4380
rect 15194 4378 15200 4380
rect 14954 4326 14956 4378
rect 15136 4326 15138 4378
rect 14892 4324 14898 4326
rect 14954 4324 14978 4326
rect 15034 4324 15058 4326
rect 15114 4324 15138 4326
rect 15194 4324 15200 4326
rect 14892 4315 15200 4324
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 14232 3836 14540 3845
rect 14232 3834 14238 3836
rect 14294 3834 14318 3836
rect 14374 3834 14398 3836
rect 14454 3834 14478 3836
rect 14534 3834 14540 3836
rect 14294 3782 14296 3834
rect 14476 3782 14478 3834
rect 14232 3780 14238 3782
rect 14294 3780 14318 3782
rect 14374 3780 14398 3782
rect 14454 3780 14478 3782
rect 14534 3780 14540 3782
rect 14232 3771 14540 3780
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13832 2990 13860 3470
rect 14892 3292 15200 3301
rect 14892 3290 14898 3292
rect 14954 3290 14978 3292
rect 15034 3290 15058 3292
rect 15114 3290 15138 3292
rect 15194 3290 15200 3292
rect 14954 3238 14956 3290
rect 15136 3238 15138 3290
rect 14892 3236 14898 3238
rect 14954 3236 14978 3238
rect 15034 3236 15058 3238
rect 15114 3236 15138 3238
rect 15194 3236 15200 3238
rect 14892 3227 15200 3236
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 2847 2748 3155 2757
rect 2847 2746 2853 2748
rect 2909 2746 2933 2748
rect 2989 2746 3013 2748
rect 3069 2746 3093 2748
rect 3149 2746 3155 2748
rect 2909 2694 2911 2746
rect 3091 2694 3093 2746
rect 2847 2692 2853 2694
rect 2909 2692 2933 2694
rect 2989 2692 3013 2694
rect 3069 2692 3093 2694
rect 3149 2692 3155 2694
rect 2847 2683 3155 2692
rect 4448 2746 4568 2774
rect 6642 2748 6950 2757
rect 6642 2746 6648 2748
rect 6704 2746 6728 2748
rect 6784 2746 6808 2748
rect 6864 2746 6888 2748
rect 6944 2746 6950 2748
rect 4448 2650 4476 2746
rect 6704 2694 6706 2746
rect 6886 2694 6888 2746
rect 6642 2692 6648 2694
rect 6704 2692 6728 2694
rect 6784 2692 6808 2694
rect 6864 2692 6888 2694
rect 6944 2692 6950 2694
rect 6642 2683 6950 2692
rect 10437 2748 10745 2757
rect 10437 2746 10443 2748
rect 10499 2746 10523 2748
rect 10579 2746 10603 2748
rect 10659 2746 10683 2748
rect 10739 2746 10745 2748
rect 10499 2694 10501 2746
rect 10681 2694 10683 2746
rect 10437 2692 10443 2694
rect 10499 2692 10523 2694
rect 10579 2692 10603 2694
rect 10659 2692 10683 2694
rect 10739 2692 10745 2694
rect 10437 2683 10745 2692
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 13832 2514 13860 2926
rect 14232 2748 14540 2757
rect 14232 2746 14238 2748
rect 14294 2746 14318 2748
rect 14374 2746 14398 2748
rect 14454 2746 14478 2748
rect 14534 2746 14540 2748
rect 14294 2694 14296 2746
rect 14476 2694 14478 2746
rect 14232 2692 14238 2694
rect 14294 2692 14318 2694
rect 14374 2692 14398 2694
rect 14454 2692 14478 2694
rect 14534 2692 14540 2694
rect 14232 2683 14540 2692
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 32 800 60 2382
rect 3507 2204 3815 2213
rect 3507 2202 3513 2204
rect 3569 2202 3593 2204
rect 3649 2202 3673 2204
rect 3729 2202 3753 2204
rect 3809 2202 3815 2204
rect 3569 2150 3571 2202
rect 3751 2150 3753 2202
rect 3507 2148 3513 2150
rect 3569 2148 3593 2150
rect 3649 2148 3673 2150
rect 3729 2148 3753 2150
rect 3809 2148 3815 2150
rect 3507 2139 3815 2148
rect 7302 2204 7610 2213
rect 7302 2202 7308 2204
rect 7364 2202 7388 2204
rect 7444 2202 7468 2204
rect 7524 2202 7548 2204
rect 7604 2202 7610 2204
rect 7364 2150 7366 2202
rect 7546 2150 7548 2202
rect 7302 2148 7308 2150
rect 7364 2148 7388 2150
rect 7444 2148 7468 2150
rect 7524 2148 7548 2150
rect 7604 2148 7610 2150
rect 7302 2139 7610 2148
rect 11097 2204 11405 2213
rect 11097 2202 11103 2204
rect 11159 2202 11183 2204
rect 11239 2202 11263 2204
rect 11319 2202 11343 2204
rect 11399 2202 11405 2204
rect 11159 2150 11161 2202
rect 11341 2150 11343 2202
rect 11097 2148 11103 2150
rect 11159 2148 11183 2150
rect 11239 2148 11263 2150
rect 11319 2148 11343 2150
rect 11399 2148 11405 2150
rect 11097 2139 11405 2148
rect 14108 1306 14136 2382
rect 14892 2204 15200 2213
rect 14892 2202 14898 2204
rect 14954 2202 14978 2204
rect 15034 2202 15058 2204
rect 15114 2202 15138 2204
rect 15194 2202 15200 2204
rect 14954 2150 14956 2202
rect 15136 2150 15138 2202
rect 14892 2148 14898 2150
rect 14954 2148 14978 2150
rect 15034 2148 15058 2150
rect 15114 2148 15138 2150
rect 15194 2148 15200 2150
rect 14892 2139 15200 2148
rect 14108 1278 14228 1306
rect 14200 800 14228 1278
rect 18 0 74 800
rect 14186 0 14242 800
<< via2 >>
rect 2853 16890 2909 16892
rect 2933 16890 2989 16892
rect 3013 16890 3069 16892
rect 3093 16890 3149 16892
rect 2853 16838 2899 16890
rect 2899 16838 2909 16890
rect 2933 16838 2963 16890
rect 2963 16838 2975 16890
rect 2975 16838 2989 16890
rect 3013 16838 3027 16890
rect 3027 16838 3039 16890
rect 3039 16838 3069 16890
rect 3093 16838 3103 16890
rect 3103 16838 3149 16890
rect 2853 16836 2909 16838
rect 2933 16836 2989 16838
rect 3013 16836 3069 16838
rect 3093 16836 3149 16838
rect 6648 16890 6704 16892
rect 6728 16890 6784 16892
rect 6808 16890 6864 16892
rect 6888 16890 6944 16892
rect 6648 16838 6694 16890
rect 6694 16838 6704 16890
rect 6728 16838 6758 16890
rect 6758 16838 6770 16890
rect 6770 16838 6784 16890
rect 6808 16838 6822 16890
rect 6822 16838 6834 16890
rect 6834 16838 6864 16890
rect 6888 16838 6898 16890
rect 6898 16838 6944 16890
rect 6648 16836 6704 16838
rect 6728 16836 6784 16838
rect 6808 16836 6864 16838
rect 6888 16836 6944 16838
rect 10443 16890 10499 16892
rect 10523 16890 10579 16892
rect 10603 16890 10659 16892
rect 10683 16890 10739 16892
rect 10443 16838 10489 16890
rect 10489 16838 10499 16890
rect 10523 16838 10553 16890
rect 10553 16838 10565 16890
rect 10565 16838 10579 16890
rect 10603 16838 10617 16890
rect 10617 16838 10629 16890
rect 10629 16838 10659 16890
rect 10683 16838 10693 16890
rect 10693 16838 10739 16890
rect 10443 16836 10499 16838
rect 10523 16836 10579 16838
rect 10603 16836 10659 16838
rect 10683 16836 10739 16838
rect 14238 16890 14294 16892
rect 14318 16890 14374 16892
rect 14398 16890 14454 16892
rect 14478 16890 14534 16892
rect 14238 16838 14284 16890
rect 14284 16838 14294 16890
rect 14318 16838 14348 16890
rect 14348 16838 14360 16890
rect 14360 16838 14374 16890
rect 14398 16838 14412 16890
rect 14412 16838 14424 16890
rect 14424 16838 14454 16890
rect 14478 16838 14488 16890
rect 14488 16838 14534 16890
rect 14238 16836 14294 16838
rect 14318 16836 14374 16838
rect 14398 16836 14454 16838
rect 14478 16836 14534 16838
rect 3513 16346 3569 16348
rect 3593 16346 3649 16348
rect 3673 16346 3729 16348
rect 3753 16346 3809 16348
rect 3513 16294 3559 16346
rect 3559 16294 3569 16346
rect 3593 16294 3623 16346
rect 3623 16294 3635 16346
rect 3635 16294 3649 16346
rect 3673 16294 3687 16346
rect 3687 16294 3699 16346
rect 3699 16294 3729 16346
rect 3753 16294 3763 16346
rect 3763 16294 3809 16346
rect 3513 16292 3569 16294
rect 3593 16292 3649 16294
rect 3673 16292 3729 16294
rect 3753 16292 3809 16294
rect 7308 16346 7364 16348
rect 7388 16346 7444 16348
rect 7468 16346 7524 16348
rect 7548 16346 7604 16348
rect 7308 16294 7354 16346
rect 7354 16294 7364 16346
rect 7388 16294 7418 16346
rect 7418 16294 7430 16346
rect 7430 16294 7444 16346
rect 7468 16294 7482 16346
rect 7482 16294 7494 16346
rect 7494 16294 7524 16346
rect 7548 16294 7558 16346
rect 7558 16294 7604 16346
rect 7308 16292 7364 16294
rect 7388 16292 7444 16294
rect 7468 16292 7524 16294
rect 7548 16292 7604 16294
rect 2853 15802 2909 15804
rect 2933 15802 2989 15804
rect 3013 15802 3069 15804
rect 3093 15802 3149 15804
rect 2853 15750 2899 15802
rect 2899 15750 2909 15802
rect 2933 15750 2963 15802
rect 2963 15750 2975 15802
rect 2975 15750 2989 15802
rect 3013 15750 3027 15802
rect 3027 15750 3039 15802
rect 3039 15750 3069 15802
rect 3093 15750 3103 15802
rect 3103 15750 3149 15802
rect 2853 15748 2909 15750
rect 2933 15748 2989 15750
rect 3013 15748 3069 15750
rect 3093 15748 3149 15750
rect 1490 15136 1546 15192
rect 3513 15258 3569 15260
rect 3593 15258 3649 15260
rect 3673 15258 3729 15260
rect 3753 15258 3809 15260
rect 3513 15206 3559 15258
rect 3559 15206 3569 15258
rect 3593 15206 3623 15258
rect 3623 15206 3635 15258
rect 3635 15206 3649 15258
rect 3673 15206 3687 15258
rect 3687 15206 3699 15258
rect 3699 15206 3729 15258
rect 3753 15206 3763 15258
rect 3763 15206 3809 15258
rect 3513 15204 3569 15206
rect 3593 15204 3649 15206
rect 3673 15204 3729 15206
rect 3753 15204 3809 15206
rect 2853 14714 2909 14716
rect 2933 14714 2989 14716
rect 3013 14714 3069 14716
rect 3093 14714 3149 14716
rect 2853 14662 2899 14714
rect 2899 14662 2909 14714
rect 2933 14662 2963 14714
rect 2963 14662 2975 14714
rect 2975 14662 2989 14714
rect 3013 14662 3027 14714
rect 3027 14662 3039 14714
rect 3039 14662 3069 14714
rect 3093 14662 3103 14714
rect 3103 14662 3149 14714
rect 2853 14660 2909 14662
rect 2933 14660 2989 14662
rect 3013 14660 3069 14662
rect 3093 14660 3149 14662
rect 3513 14170 3569 14172
rect 3593 14170 3649 14172
rect 3673 14170 3729 14172
rect 3753 14170 3809 14172
rect 3513 14118 3559 14170
rect 3559 14118 3569 14170
rect 3593 14118 3623 14170
rect 3623 14118 3635 14170
rect 3635 14118 3649 14170
rect 3673 14118 3687 14170
rect 3687 14118 3699 14170
rect 3699 14118 3729 14170
rect 3753 14118 3763 14170
rect 3763 14118 3809 14170
rect 3513 14116 3569 14118
rect 3593 14116 3649 14118
rect 3673 14116 3729 14118
rect 3753 14116 3809 14118
rect 2853 13626 2909 13628
rect 2933 13626 2989 13628
rect 3013 13626 3069 13628
rect 3093 13626 3149 13628
rect 2853 13574 2899 13626
rect 2899 13574 2909 13626
rect 2933 13574 2963 13626
rect 2963 13574 2975 13626
rect 2975 13574 2989 13626
rect 3013 13574 3027 13626
rect 3027 13574 3039 13626
rect 3039 13574 3069 13626
rect 3093 13574 3103 13626
rect 3103 13574 3149 13626
rect 2853 13572 2909 13574
rect 2933 13572 2989 13574
rect 3013 13572 3069 13574
rect 3093 13572 3149 13574
rect 3513 13082 3569 13084
rect 3593 13082 3649 13084
rect 3673 13082 3729 13084
rect 3753 13082 3809 13084
rect 3513 13030 3559 13082
rect 3559 13030 3569 13082
rect 3593 13030 3623 13082
rect 3623 13030 3635 13082
rect 3635 13030 3649 13082
rect 3673 13030 3687 13082
rect 3687 13030 3699 13082
rect 3699 13030 3729 13082
rect 3753 13030 3763 13082
rect 3763 13030 3809 13082
rect 3513 13028 3569 13030
rect 3593 13028 3649 13030
rect 3673 13028 3729 13030
rect 3753 13028 3809 13030
rect 2853 12538 2909 12540
rect 2933 12538 2989 12540
rect 3013 12538 3069 12540
rect 3093 12538 3149 12540
rect 2853 12486 2899 12538
rect 2899 12486 2909 12538
rect 2933 12486 2963 12538
rect 2963 12486 2975 12538
rect 2975 12486 2989 12538
rect 3013 12486 3027 12538
rect 3027 12486 3039 12538
rect 3039 12486 3069 12538
rect 3093 12486 3103 12538
rect 3103 12486 3149 12538
rect 2853 12484 2909 12486
rect 2933 12484 2989 12486
rect 3013 12484 3069 12486
rect 3093 12484 3149 12486
rect 6648 15802 6704 15804
rect 6728 15802 6784 15804
rect 6808 15802 6864 15804
rect 6888 15802 6944 15804
rect 6648 15750 6694 15802
rect 6694 15750 6704 15802
rect 6728 15750 6758 15802
rect 6758 15750 6770 15802
rect 6770 15750 6784 15802
rect 6808 15750 6822 15802
rect 6822 15750 6834 15802
rect 6834 15750 6864 15802
rect 6888 15750 6898 15802
rect 6898 15750 6944 15802
rect 6648 15748 6704 15750
rect 6728 15748 6784 15750
rect 6808 15748 6864 15750
rect 6888 15748 6944 15750
rect 6648 14714 6704 14716
rect 6728 14714 6784 14716
rect 6808 14714 6864 14716
rect 6888 14714 6944 14716
rect 6648 14662 6694 14714
rect 6694 14662 6704 14714
rect 6728 14662 6758 14714
rect 6758 14662 6770 14714
rect 6770 14662 6784 14714
rect 6808 14662 6822 14714
rect 6822 14662 6834 14714
rect 6834 14662 6864 14714
rect 6888 14662 6898 14714
rect 6898 14662 6944 14714
rect 6648 14660 6704 14662
rect 6728 14660 6784 14662
rect 6808 14660 6864 14662
rect 6888 14660 6944 14662
rect 7308 15258 7364 15260
rect 7388 15258 7444 15260
rect 7468 15258 7524 15260
rect 7548 15258 7604 15260
rect 7308 15206 7354 15258
rect 7354 15206 7364 15258
rect 7388 15206 7418 15258
rect 7418 15206 7430 15258
rect 7430 15206 7444 15258
rect 7468 15206 7482 15258
rect 7482 15206 7494 15258
rect 7494 15206 7524 15258
rect 7548 15206 7558 15258
rect 7558 15206 7604 15258
rect 7308 15204 7364 15206
rect 7388 15204 7444 15206
rect 7468 15204 7524 15206
rect 7548 15204 7604 15206
rect 6648 13626 6704 13628
rect 6728 13626 6784 13628
rect 6808 13626 6864 13628
rect 6888 13626 6944 13628
rect 6648 13574 6694 13626
rect 6694 13574 6704 13626
rect 6728 13574 6758 13626
rect 6758 13574 6770 13626
rect 6770 13574 6784 13626
rect 6808 13574 6822 13626
rect 6822 13574 6834 13626
rect 6834 13574 6864 13626
rect 6888 13574 6898 13626
rect 6898 13574 6944 13626
rect 6648 13572 6704 13574
rect 6728 13572 6784 13574
rect 6808 13572 6864 13574
rect 6888 13572 6944 13574
rect 2853 11450 2909 11452
rect 2933 11450 2989 11452
rect 3013 11450 3069 11452
rect 3093 11450 3149 11452
rect 2853 11398 2899 11450
rect 2899 11398 2909 11450
rect 2933 11398 2963 11450
rect 2963 11398 2975 11450
rect 2975 11398 2989 11450
rect 3013 11398 3027 11450
rect 3027 11398 3039 11450
rect 3039 11398 3069 11450
rect 3093 11398 3103 11450
rect 3103 11398 3149 11450
rect 2853 11396 2909 11398
rect 2933 11396 2989 11398
rect 3013 11396 3069 11398
rect 3093 11396 3149 11398
rect 3513 11994 3569 11996
rect 3593 11994 3649 11996
rect 3673 11994 3729 11996
rect 3753 11994 3809 11996
rect 3513 11942 3559 11994
rect 3559 11942 3569 11994
rect 3593 11942 3623 11994
rect 3623 11942 3635 11994
rect 3635 11942 3649 11994
rect 3673 11942 3687 11994
rect 3687 11942 3699 11994
rect 3699 11942 3729 11994
rect 3753 11942 3763 11994
rect 3763 11942 3809 11994
rect 3513 11940 3569 11942
rect 3593 11940 3649 11942
rect 3673 11940 3729 11942
rect 3753 11940 3809 11942
rect 6648 12538 6704 12540
rect 6728 12538 6784 12540
rect 6808 12538 6864 12540
rect 6888 12538 6944 12540
rect 6648 12486 6694 12538
rect 6694 12486 6704 12538
rect 6728 12486 6758 12538
rect 6758 12486 6770 12538
rect 6770 12486 6784 12538
rect 6808 12486 6822 12538
rect 6822 12486 6834 12538
rect 6834 12486 6864 12538
rect 6888 12486 6898 12538
rect 6898 12486 6944 12538
rect 6648 12484 6704 12486
rect 6728 12484 6784 12486
rect 6808 12484 6864 12486
rect 6888 12484 6944 12486
rect 7308 14170 7364 14172
rect 7388 14170 7444 14172
rect 7468 14170 7524 14172
rect 7548 14170 7604 14172
rect 7308 14118 7354 14170
rect 7354 14118 7364 14170
rect 7388 14118 7418 14170
rect 7418 14118 7430 14170
rect 7430 14118 7444 14170
rect 7468 14118 7482 14170
rect 7482 14118 7494 14170
rect 7494 14118 7524 14170
rect 7548 14118 7558 14170
rect 7558 14118 7604 14170
rect 7308 14116 7364 14118
rect 7388 14116 7444 14118
rect 7468 14116 7524 14118
rect 7548 14116 7604 14118
rect 11103 16346 11159 16348
rect 11183 16346 11239 16348
rect 11263 16346 11319 16348
rect 11343 16346 11399 16348
rect 11103 16294 11149 16346
rect 11149 16294 11159 16346
rect 11183 16294 11213 16346
rect 11213 16294 11225 16346
rect 11225 16294 11239 16346
rect 11263 16294 11277 16346
rect 11277 16294 11289 16346
rect 11289 16294 11319 16346
rect 11343 16294 11353 16346
rect 11353 16294 11399 16346
rect 11103 16292 11159 16294
rect 11183 16292 11239 16294
rect 11263 16292 11319 16294
rect 11343 16292 11399 16294
rect 14898 16346 14954 16348
rect 14978 16346 15034 16348
rect 15058 16346 15114 16348
rect 15138 16346 15194 16348
rect 14898 16294 14944 16346
rect 14944 16294 14954 16346
rect 14978 16294 15008 16346
rect 15008 16294 15020 16346
rect 15020 16294 15034 16346
rect 15058 16294 15072 16346
rect 15072 16294 15084 16346
rect 15084 16294 15114 16346
rect 15138 16294 15148 16346
rect 15148 16294 15194 16346
rect 14898 16292 14954 16294
rect 14978 16292 15034 16294
rect 15058 16292 15114 16294
rect 15138 16292 15194 16294
rect 10443 15802 10499 15804
rect 10523 15802 10579 15804
rect 10603 15802 10659 15804
rect 10683 15802 10739 15804
rect 10443 15750 10489 15802
rect 10489 15750 10499 15802
rect 10523 15750 10553 15802
rect 10553 15750 10565 15802
rect 10565 15750 10579 15802
rect 10603 15750 10617 15802
rect 10617 15750 10629 15802
rect 10629 15750 10659 15802
rect 10683 15750 10693 15802
rect 10693 15750 10739 15802
rect 10443 15748 10499 15750
rect 10523 15748 10579 15750
rect 10603 15748 10659 15750
rect 10683 15748 10739 15750
rect 10443 14714 10499 14716
rect 10523 14714 10579 14716
rect 10603 14714 10659 14716
rect 10683 14714 10739 14716
rect 10443 14662 10489 14714
rect 10489 14662 10499 14714
rect 10523 14662 10553 14714
rect 10553 14662 10565 14714
rect 10565 14662 10579 14714
rect 10603 14662 10617 14714
rect 10617 14662 10629 14714
rect 10629 14662 10659 14714
rect 10683 14662 10693 14714
rect 10693 14662 10739 14714
rect 10443 14660 10499 14662
rect 10523 14660 10579 14662
rect 10603 14660 10659 14662
rect 10683 14660 10739 14662
rect 7308 13082 7364 13084
rect 7388 13082 7444 13084
rect 7468 13082 7524 13084
rect 7548 13082 7604 13084
rect 7308 13030 7354 13082
rect 7354 13030 7364 13082
rect 7388 13030 7418 13082
rect 7418 13030 7430 13082
rect 7430 13030 7444 13082
rect 7468 13030 7482 13082
rect 7482 13030 7494 13082
rect 7494 13030 7524 13082
rect 7548 13030 7558 13082
rect 7558 13030 7604 13082
rect 7308 13028 7364 13030
rect 7388 13028 7444 13030
rect 7468 13028 7524 13030
rect 7548 13028 7604 13030
rect 6648 11450 6704 11452
rect 6728 11450 6784 11452
rect 6808 11450 6864 11452
rect 6888 11450 6944 11452
rect 6648 11398 6694 11450
rect 6694 11398 6704 11450
rect 6728 11398 6758 11450
rect 6758 11398 6770 11450
rect 6770 11398 6784 11450
rect 6808 11398 6822 11450
rect 6822 11398 6834 11450
rect 6834 11398 6864 11450
rect 6888 11398 6898 11450
rect 6898 11398 6944 11450
rect 6648 11396 6704 11398
rect 6728 11396 6784 11398
rect 6808 11396 6864 11398
rect 6888 11396 6944 11398
rect 3513 10906 3569 10908
rect 3593 10906 3649 10908
rect 3673 10906 3729 10908
rect 3753 10906 3809 10908
rect 3513 10854 3559 10906
rect 3559 10854 3569 10906
rect 3593 10854 3623 10906
rect 3623 10854 3635 10906
rect 3635 10854 3649 10906
rect 3673 10854 3687 10906
rect 3687 10854 3699 10906
rect 3699 10854 3729 10906
rect 3753 10854 3763 10906
rect 3763 10854 3809 10906
rect 3513 10852 3569 10854
rect 3593 10852 3649 10854
rect 3673 10852 3729 10854
rect 3753 10852 3809 10854
rect 2853 10362 2909 10364
rect 2933 10362 2989 10364
rect 3013 10362 3069 10364
rect 3093 10362 3149 10364
rect 2853 10310 2899 10362
rect 2899 10310 2909 10362
rect 2933 10310 2963 10362
rect 2963 10310 2975 10362
rect 2975 10310 2989 10362
rect 3013 10310 3027 10362
rect 3027 10310 3039 10362
rect 3039 10310 3069 10362
rect 3093 10310 3103 10362
rect 3103 10310 3149 10362
rect 2853 10308 2909 10310
rect 2933 10308 2989 10310
rect 3013 10308 3069 10310
rect 3093 10308 3149 10310
rect 2853 9274 2909 9276
rect 2933 9274 2989 9276
rect 3013 9274 3069 9276
rect 3093 9274 3149 9276
rect 2853 9222 2899 9274
rect 2899 9222 2909 9274
rect 2933 9222 2963 9274
rect 2963 9222 2975 9274
rect 2975 9222 2989 9274
rect 3013 9222 3027 9274
rect 3027 9222 3039 9274
rect 3039 9222 3069 9274
rect 3093 9222 3103 9274
rect 3103 9222 3149 9274
rect 2853 9220 2909 9222
rect 2933 9220 2989 9222
rect 3013 9220 3069 9222
rect 3093 9220 3149 9222
rect 2853 8186 2909 8188
rect 2933 8186 2989 8188
rect 3013 8186 3069 8188
rect 3093 8186 3149 8188
rect 2853 8134 2899 8186
rect 2899 8134 2909 8186
rect 2933 8134 2963 8186
rect 2963 8134 2975 8186
rect 2975 8134 2989 8186
rect 3013 8134 3027 8186
rect 3027 8134 3039 8186
rect 3039 8134 3069 8186
rect 3093 8134 3103 8186
rect 3103 8134 3149 8186
rect 2853 8132 2909 8134
rect 2933 8132 2989 8134
rect 3013 8132 3069 8134
rect 3093 8132 3149 8134
rect 3513 9818 3569 9820
rect 3593 9818 3649 9820
rect 3673 9818 3729 9820
rect 3753 9818 3809 9820
rect 3513 9766 3559 9818
rect 3559 9766 3569 9818
rect 3593 9766 3623 9818
rect 3623 9766 3635 9818
rect 3635 9766 3649 9818
rect 3673 9766 3687 9818
rect 3687 9766 3699 9818
rect 3699 9766 3729 9818
rect 3753 9766 3763 9818
rect 3763 9766 3809 9818
rect 3513 9764 3569 9766
rect 3593 9764 3649 9766
rect 3673 9764 3729 9766
rect 3753 9764 3809 9766
rect 3513 8730 3569 8732
rect 3593 8730 3649 8732
rect 3673 8730 3729 8732
rect 3753 8730 3809 8732
rect 3513 8678 3559 8730
rect 3559 8678 3569 8730
rect 3593 8678 3623 8730
rect 3623 8678 3635 8730
rect 3635 8678 3649 8730
rect 3673 8678 3687 8730
rect 3687 8678 3699 8730
rect 3699 8678 3729 8730
rect 3753 8678 3763 8730
rect 3763 8678 3809 8730
rect 3513 8676 3569 8678
rect 3593 8676 3649 8678
rect 3673 8676 3729 8678
rect 3753 8676 3809 8678
rect 3513 7642 3569 7644
rect 3593 7642 3649 7644
rect 3673 7642 3729 7644
rect 3753 7642 3809 7644
rect 3513 7590 3559 7642
rect 3559 7590 3569 7642
rect 3593 7590 3623 7642
rect 3623 7590 3635 7642
rect 3635 7590 3649 7642
rect 3673 7590 3687 7642
rect 3687 7590 3699 7642
rect 3699 7590 3729 7642
rect 3753 7590 3763 7642
rect 3763 7590 3809 7642
rect 3513 7588 3569 7590
rect 3593 7588 3649 7590
rect 3673 7588 3729 7590
rect 3753 7588 3809 7590
rect 2853 7098 2909 7100
rect 2933 7098 2989 7100
rect 3013 7098 3069 7100
rect 3093 7098 3149 7100
rect 2853 7046 2899 7098
rect 2899 7046 2909 7098
rect 2933 7046 2963 7098
rect 2963 7046 2975 7098
rect 2975 7046 2989 7098
rect 3013 7046 3027 7098
rect 3027 7046 3039 7098
rect 3039 7046 3069 7098
rect 3093 7046 3103 7098
rect 3103 7046 3149 7098
rect 2853 7044 2909 7046
rect 2933 7044 2989 7046
rect 3013 7044 3069 7046
rect 3093 7044 3149 7046
rect 2853 6010 2909 6012
rect 2933 6010 2989 6012
rect 3013 6010 3069 6012
rect 3093 6010 3149 6012
rect 2853 5958 2899 6010
rect 2899 5958 2909 6010
rect 2933 5958 2963 6010
rect 2963 5958 2975 6010
rect 2975 5958 2989 6010
rect 3013 5958 3027 6010
rect 3027 5958 3039 6010
rect 3039 5958 3069 6010
rect 3093 5958 3103 6010
rect 3103 5958 3149 6010
rect 2853 5956 2909 5958
rect 2933 5956 2989 5958
rect 3013 5956 3069 5958
rect 3093 5956 3149 5958
rect 2853 4922 2909 4924
rect 2933 4922 2989 4924
rect 3013 4922 3069 4924
rect 3093 4922 3149 4924
rect 2853 4870 2899 4922
rect 2899 4870 2909 4922
rect 2933 4870 2963 4922
rect 2963 4870 2975 4922
rect 2975 4870 2989 4922
rect 3013 4870 3027 4922
rect 3027 4870 3039 4922
rect 3039 4870 3069 4922
rect 3093 4870 3103 4922
rect 3103 4870 3149 4922
rect 2853 4868 2909 4870
rect 2933 4868 2989 4870
rect 3013 4868 3069 4870
rect 3093 4868 3149 4870
rect 3513 6554 3569 6556
rect 3593 6554 3649 6556
rect 3673 6554 3729 6556
rect 3753 6554 3809 6556
rect 3513 6502 3559 6554
rect 3559 6502 3569 6554
rect 3593 6502 3623 6554
rect 3623 6502 3635 6554
rect 3635 6502 3649 6554
rect 3673 6502 3687 6554
rect 3687 6502 3699 6554
rect 3699 6502 3729 6554
rect 3753 6502 3763 6554
rect 3763 6502 3809 6554
rect 3513 6500 3569 6502
rect 3593 6500 3649 6502
rect 3673 6500 3729 6502
rect 3753 6500 3809 6502
rect 3513 5466 3569 5468
rect 3593 5466 3649 5468
rect 3673 5466 3729 5468
rect 3753 5466 3809 5468
rect 3513 5414 3559 5466
rect 3559 5414 3569 5466
rect 3593 5414 3623 5466
rect 3623 5414 3635 5466
rect 3635 5414 3649 5466
rect 3673 5414 3687 5466
rect 3687 5414 3699 5466
rect 3699 5414 3729 5466
rect 3753 5414 3763 5466
rect 3763 5414 3809 5466
rect 3513 5412 3569 5414
rect 3593 5412 3649 5414
rect 3673 5412 3729 5414
rect 3753 5412 3809 5414
rect 3513 4378 3569 4380
rect 3593 4378 3649 4380
rect 3673 4378 3729 4380
rect 3753 4378 3809 4380
rect 3513 4326 3559 4378
rect 3559 4326 3569 4378
rect 3593 4326 3623 4378
rect 3623 4326 3635 4378
rect 3635 4326 3649 4378
rect 3673 4326 3687 4378
rect 3687 4326 3699 4378
rect 3699 4326 3729 4378
rect 3753 4326 3763 4378
rect 3763 4326 3809 4378
rect 3513 4324 3569 4326
rect 3593 4324 3649 4326
rect 3673 4324 3729 4326
rect 3753 4324 3809 4326
rect 2853 3834 2909 3836
rect 2933 3834 2989 3836
rect 3013 3834 3069 3836
rect 3093 3834 3149 3836
rect 2853 3782 2899 3834
rect 2899 3782 2909 3834
rect 2933 3782 2963 3834
rect 2963 3782 2975 3834
rect 2975 3782 2989 3834
rect 3013 3782 3027 3834
rect 3027 3782 3039 3834
rect 3039 3782 3069 3834
rect 3093 3782 3103 3834
rect 3103 3782 3149 3834
rect 2853 3780 2909 3782
rect 2933 3780 2989 3782
rect 3013 3780 3069 3782
rect 3093 3780 3149 3782
rect 6648 10362 6704 10364
rect 6728 10362 6784 10364
rect 6808 10362 6864 10364
rect 6888 10362 6944 10364
rect 6648 10310 6694 10362
rect 6694 10310 6704 10362
rect 6728 10310 6758 10362
rect 6758 10310 6770 10362
rect 6770 10310 6784 10362
rect 6808 10310 6822 10362
rect 6822 10310 6834 10362
rect 6834 10310 6864 10362
rect 6888 10310 6898 10362
rect 6898 10310 6944 10362
rect 6648 10308 6704 10310
rect 6728 10308 6784 10310
rect 6808 10308 6864 10310
rect 6888 10308 6944 10310
rect 5446 9016 5502 9072
rect 7308 11994 7364 11996
rect 7388 11994 7444 11996
rect 7468 11994 7524 11996
rect 7548 11994 7604 11996
rect 7308 11942 7354 11994
rect 7354 11942 7364 11994
rect 7388 11942 7418 11994
rect 7418 11942 7430 11994
rect 7430 11942 7444 11994
rect 7468 11942 7482 11994
rect 7482 11942 7494 11994
rect 7494 11942 7524 11994
rect 7548 11942 7558 11994
rect 7558 11942 7604 11994
rect 7308 11940 7364 11942
rect 7388 11940 7444 11942
rect 7468 11940 7524 11942
rect 7548 11940 7604 11942
rect 7308 10906 7364 10908
rect 7388 10906 7444 10908
rect 7468 10906 7524 10908
rect 7548 10906 7604 10908
rect 7308 10854 7354 10906
rect 7354 10854 7364 10906
rect 7388 10854 7418 10906
rect 7418 10854 7430 10906
rect 7430 10854 7444 10906
rect 7468 10854 7482 10906
rect 7482 10854 7494 10906
rect 7494 10854 7524 10906
rect 7548 10854 7558 10906
rect 7558 10854 7604 10906
rect 7308 10852 7364 10854
rect 7388 10852 7444 10854
rect 7468 10852 7524 10854
rect 7548 10852 7604 10854
rect 7308 9818 7364 9820
rect 7388 9818 7444 9820
rect 7468 9818 7524 9820
rect 7548 9818 7604 9820
rect 7308 9766 7354 9818
rect 7354 9766 7364 9818
rect 7388 9766 7418 9818
rect 7418 9766 7430 9818
rect 7430 9766 7444 9818
rect 7468 9766 7482 9818
rect 7482 9766 7494 9818
rect 7494 9766 7524 9818
rect 7548 9766 7558 9818
rect 7558 9766 7604 9818
rect 7308 9764 7364 9766
rect 7388 9764 7444 9766
rect 7468 9764 7524 9766
rect 7548 9764 7604 9766
rect 6648 9274 6704 9276
rect 6728 9274 6784 9276
rect 6808 9274 6864 9276
rect 6888 9274 6944 9276
rect 6648 9222 6694 9274
rect 6694 9222 6704 9274
rect 6728 9222 6758 9274
rect 6758 9222 6770 9274
rect 6770 9222 6784 9274
rect 6808 9222 6822 9274
rect 6822 9222 6834 9274
rect 6834 9222 6864 9274
rect 6888 9222 6898 9274
rect 6898 9222 6944 9274
rect 6648 9220 6704 9222
rect 6728 9220 6784 9222
rect 6808 9220 6864 9222
rect 6888 9220 6944 9222
rect 3513 3290 3569 3292
rect 3593 3290 3649 3292
rect 3673 3290 3729 3292
rect 3753 3290 3809 3292
rect 3513 3238 3559 3290
rect 3559 3238 3569 3290
rect 3593 3238 3623 3290
rect 3623 3238 3635 3290
rect 3635 3238 3649 3290
rect 3673 3238 3687 3290
rect 3687 3238 3699 3290
rect 3699 3238 3729 3290
rect 3753 3238 3763 3290
rect 3763 3238 3809 3290
rect 3513 3236 3569 3238
rect 3593 3236 3649 3238
rect 3673 3236 3729 3238
rect 3753 3236 3809 3238
rect 6648 8186 6704 8188
rect 6728 8186 6784 8188
rect 6808 8186 6864 8188
rect 6888 8186 6944 8188
rect 6648 8134 6694 8186
rect 6694 8134 6704 8186
rect 6728 8134 6758 8186
rect 6758 8134 6770 8186
rect 6770 8134 6784 8186
rect 6808 8134 6822 8186
rect 6822 8134 6834 8186
rect 6834 8134 6864 8186
rect 6888 8134 6898 8186
rect 6898 8134 6944 8186
rect 6648 8132 6704 8134
rect 6728 8132 6784 8134
rect 6808 8132 6864 8134
rect 6888 8132 6944 8134
rect 7308 8730 7364 8732
rect 7388 8730 7444 8732
rect 7468 8730 7524 8732
rect 7548 8730 7604 8732
rect 7308 8678 7354 8730
rect 7354 8678 7364 8730
rect 7388 8678 7418 8730
rect 7418 8678 7430 8730
rect 7430 8678 7444 8730
rect 7468 8678 7482 8730
rect 7482 8678 7494 8730
rect 7494 8678 7524 8730
rect 7548 8678 7558 8730
rect 7558 8678 7604 8730
rect 7308 8676 7364 8678
rect 7388 8676 7444 8678
rect 7468 8676 7524 8678
rect 7548 8676 7604 8678
rect 7308 7642 7364 7644
rect 7388 7642 7444 7644
rect 7468 7642 7524 7644
rect 7548 7642 7604 7644
rect 7308 7590 7354 7642
rect 7354 7590 7364 7642
rect 7388 7590 7418 7642
rect 7418 7590 7430 7642
rect 7430 7590 7444 7642
rect 7468 7590 7482 7642
rect 7482 7590 7494 7642
rect 7494 7590 7524 7642
rect 7548 7590 7558 7642
rect 7558 7590 7604 7642
rect 7308 7588 7364 7590
rect 7388 7588 7444 7590
rect 7468 7588 7524 7590
rect 7548 7588 7604 7590
rect 9586 9036 9642 9072
rect 9586 9016 9588 9036
rect 9588 9016 9640 9036
rect 9640 9016 9642 9036
rect 6648 7098 6704 7100
rect 6728 7098 6784 7100
rect 6808 7098 6864 7100
rect 6888 7098 6944 7100
rect 6648 7046 6694 7098
rect 6694 7046 6704 7098
rect 6728 7046 6758 7098
rect 6758 7046 6770 7098
rect 6770 7046 6784 7098
rect 6808 7046 6822 7098
rect 6822 7046 6834 7098
rect 6834 7046 6864 7098
rect 6888 7046 6898 7098
rect 6898 7046 6944 7098
rect 6648 7044 6704 7046
rect 6728 7044 6784 7046
rect 6808 7044 6864 7046
rect 6888 7044 6944 7046
rect 6648 6010 6704 6012
rect 6728 6010 6784 6012
rect 6808 6010 6864 6012
rect 6888 6010 6944 6012
rect 6648 5958 6694 6010
rect 6694 5958 6704 6010
rect 6728 5958 6758 6010
rect 6758 5958 6770 6010
rect 6770 5958 6784 6010
rect 6808 5958 6822 6010
rect 6822 5958 6834 6010
rect 6834 5958 6864 6010
rect 6888 5958 6898 6010
rect 6898 5958 6944 6010
rect 6648 5956 6704 5958
rect 6728 5956 6784 5958
rect 6808 5956 6864 5958
rect 6888 5956 6944 5958
rect 7308 6554 7364 6556
rect 7388 6554 7444 6556
rect 7468 6554 7524 6556
rect 7548 6554 7604 6556
rect 7308 6502 7354 6554
rect 7354 6502 7364 6554
rect 7388 6502 7418 6554
rect 7418 6502 7430 6554
rect 7430 6502 7444 6554
rect 7468 6502 7482 6554
rect 7482 6502 7494 6554
rect 7494 6502 7524 6554
rect 7548 6502 7558 6554
rect 7558 6502 7604 6554
rect 7308 6500 7364 6502
rect 7388 6500 7444 6502
rect 7468 6500 7524 6502
rect 7548 6500 7604 6502
rect 11103 15258 11159 15260
rect 11183 15258 11239 15260
rect 11263 15258 11319 15260
rect 11343 15258 11399 15260
rect 11103 15206 11149 15258
rect 11149 15206 11159 15258
rect 11183 15206 11213 15258
rect 11213 15206 11225 15258
rect 11225 15206 11239 15258
rect 11263 15206 11277 15258
rect 11277 15206 11289 15258
rect 11289 15206 11319 15258
rect 11343 15206 11353 15258
rect 11353 15206 11399 15258
rect 11103 15204 11159 15206
rect 11183 15204 11239 15206
rect 11263 15204 11319 15206
rect 11343 15204 11399 15206
rect 14238 15802 14294 15804
rect 14318 15802 14374 15804
rect 14398 15802 14454 15804
rect 14478 15802 14534 15804
rect 14238 15750 14284 15802
rect 14284 15750 14294 15802
rect 14318 15750 14348 15802
rect 14348 15750 14360 15802
rect 14360 15750 14374 15802
rect 14398 15750 14412 15802
rect 14412 15750 14424 15802
rect 14424 15750 14454 15802
rect 14478 15750 14488 15802
rect 14488 15750 14534 15802
rect 14238 15748 14294 15750
rect 14318 15748 14374 15750
rect 14398 15748 14454 15750
rect 14478 15748 14534 15750
rect 11103 14170 11159 14172
rect 11183 14170 11239 14172
rect 11263 14170 11319 14172
rect 11343 14170 11399 14172
rect 11103 14118 11149 14170
rect 11149 14118 11159 14170
rect 11183 14118 11213 14170
rect 11213 14118 11225 14170
rect 11225 14118 11239 14170
rect 11263 14118 11277 14170
rect 11277 14118 11289 14170
rect 11289 14118 11319 14170
rect 11343 14118 11353 14170
rect 11353 14118 11399 14170
rect 11103 14116 11159 14118
rect 11183 14116 11239 14118
rect 11263 14116 11319 14118
rect 11343 14116 11399 14118
rect 10443 13626 10499 13628
rect 10523 13626 10579 13628
rect 10603 13626 10659 13628
rect 10683 13626 10739 13628
rect 10443 13574 10489 13626
rect 10489 13574 10499 13626
rect 10523 13574 10553 13626
rect 10553 13574 10565 13626
rect 10565 13574 10579 13626
rect 10603 13574 10617 13626
rect 10617 13574 10629 13626
rect 10629 13574 10659 13626
rect 10683 13574 10693 13626
rect 10693 13574 10739 13626
rect 10443 13572 10499 13574
rect 10523 13572 10579 13574
rect 10603 13572 10659 13574
rect 10683 13572 10739 13574
rect 11103 13082 11159 13084
rect 11183 13082 11239 13084
rect 11263 13082 11319 13084
rect 11343 13082 11399 13084
rect 11103 13030 11149 13082
rect 11149 13030 11159 13082
rect 11183 13030 11213 13082
rect 11213 13030 11225 13082
rect 11225 13030 11239 13082
rect 11263 13030 11277 13082
rect 11277 13030 11289 13082
rect 11289 13030 11319 13082
rect 11343 13030 11353 13082
rect 11353 13030 11399 13082
rect 11103 13028 11159 13030
rect 11183 13028 11239 13030
rect 11263 13028 11319 13030
rect 11343 13028 11399 13030
rect 10443 12538 10499 12540
rect 10523 12538 10579 12540
rect 10603 12538 10659 12540
rect 10683 12538 10739 12540
rect 10443 12486 10489 12538
rect 10489 12486 10499 12538
rect 10523 12486 10553 12538
rect 10553 12486 10565 12538
rect 10565 12486 10579 12538
rect 10603 12486 10617 12538
rect 10617 12486 10629 12538
rect 10629 12486 10659 12538
rect 10683 12486 10693 12538
rect 10693 12486 10739 12538
rect 10443 12484 10499 12486
rect 10523 12484 10579 12486
rect 10603 12484 10659 12486
rect 10683 12484 10739 12486
rect 11103 11994 11159 11996
rect 11183 11994 11239 11996
rect 11263 11994 11319 11996
rect 11343 11994 11399 11996
rect 11103 11942 11149 11994
rect 11149 11942 11159 11994
rect 11183 11942 11213 11994
rect 11213 11942 11225 11994
rect 11225 11942 11239 11994
rect 11263 11942 11277 11994
rect 11277 11942 11289 11994
rect 11289 11942 11319 11994
rect 11343 11942 11353 11994
rect 11353 11942 11399 11994
rect 11103 11940 11159 11942
rect 11183 11940 11239 11942
rect 11263 11940 11319 11942
rect 11343 11940 11399 11942
rect 10443 11450 10499 11452
rect 10523 11450 10579 11452
rect 10603 11450 10659 11452
rect 10683 11450 10739 11452
rect 10443 11398 10489 11450
rect 10489 11398 10499 11450
rect 10523 11398 10553 11450
rect 10553 11398 10565 11450
rect 10565 11398 10579 11450
rect 10603 11398 10617 11450
rect 10617 11398 10629 11450
rect 10629 11398 10659 11450
rect 10683 11398 10693 11450
rect 10693 11398 10739 11450
rect 10443 11396 10499 11398
rect 10523 11396 10579 11398
rect 10603 11396 10659 11398
rect 10683 11396 10739 11398
rect 10443 10362 10499 10364
rect 10523 10362 10579 10364
rect 10603 10362 10659 10364
rect 10683 10362 10739 10364
rect 10443 10310 10489 10362
rect 10489 10310 10499 10362
rect 10523 10310 10553 10362
rect 10553 10310 10565 10362
rect 10565 10310 10579 10362
rect 10603 10310 10617 10362
rect 10617 10310 10629 10362
rect 10629 10310 10659 10362
rect 10683 10310 10693 10362
rect 10693 10310 10739 10362
rect 10443 10308 10499 10310
rect 10523 10308 10579 10310
rect 10603 10308 10659 10310
rect 10683 10308 10739 10310
rect 11103 10906 11159 10908
rect 11183 10906 11239 10908
rect 11263 10906 11319 10908
rect 11343 10906 11399 10908
rect 11103 10854 11149 10906
rect 11149 10854 11159 10906
rect 11183 10854 11213 10906
rect 11213 10854 11225 10906
rect 11225 10854 11239 10906
rect 11263 10854 11277 10906
rect 11277 10854 11289 10906
rect 11289 10854 11319 10906
rect 11343 10854 11353 10906
rect 11353 10854 11399 10906
rect 11103 10852 11159 10854
rect 11183 10852 11239 10854
rect 11263 10852 11319 10854
rect 11343 10852 11399 10854
rect 11103 9818 11159 9820
rect 11183 9818 11239 9820
rect 11263 9818 11319 9820
rect 11343 9818 11399 9820
rect 11103 9766 11149 9818
rect 11149 9766 11159 9818
rect 11183 9766 11213 9818
rect 11213 9766 11225 9818
rect 11225 9766 11239 9818
rect 11263 9766 11277 9818
rect 11277 9766 11289 9818
rect 11289 9766 11319 9818
rect 11343 9766 11353 9818
rect 11353 9766 11399 9818
rect 11103 9764 11159 9766
rect 11183 9764 11239 9766
rect 11263 9764 11319 9766
rect 11343 9764 11399 9766
rect 6648 4922 6704 4924
rect 6728 4922 6784 4924
rect 6808 4922 6864 4924
rect 6888 4922 6944 4924
rect 6648 4870 6694 4922
rect 6694 4870 6704 4922
rect 6728 4870 6758 4922
rect 6758 4870 6770 4922
rect 6770 4870 6784 4922
rect 6808 4870 6822 4922
rect 6822 4870 6834 4922
rect 6834 4870 6864 4922
rect 6888 4870 6898 4922
rect 6898 4870 6944 4922
rect 6648 4868 6704 4870
rect 6728 4868 6784 4870
rect 6808 4868 6864 4870
rect 6888 4868 6944 4870
rect 7308 5466 7364 5468
rect 7388 5466 7444 5468
rect 7468 5466 7524 5468
rect 7548 5466 7604 5468
rect 7308 5414 7354 5466
rect 7354 5414 7364 5466
rect 7388 5414 7418 5466
rect 7418 5414 7430 5466
rect 7430 5414 7444 5466
rect 7468 5414 7482 5466
rect 7482 5414 7494 5466
rect 7494 5414 7524 5466
rect 7548 5414 7558 5466
rect 7558 5414 7604 5466
rect 7308 5412 7364 5414
rect 7388 5412 7444 5414
rect 7468 5412 7524 5414
rect 7548 5412 7604 5414
rect 7308 4378 7364 4380
rect 7388 4378 7444 4380
rect 7468 4378 7524 4380
rect 7548 4378 7604 4380
rect 7308 4326 7354 4378
rect 7354 4326 7364 4378
rect 7388 4326 7418 4378
rect 7418 4326 7430 4378
rect 7430 4326 7444 4378
rect 7468 4326 7482 4378
rect 7482 4326 7494 4378
rect 7494 4326 7524 4378
rect 7548 4326 7558 4378
rect 7558 4326 7604 4378
rect 7308 4324 7364 4326
rect 7388 4324 7444 4326
rect 7468 4324 7524 4326
rect 7548 4324 7604 4326
rect 6648 3834 6704 3836
rect 6728 3834 6784 3836
rect 6808 3834 6864 3836
rect 6888 3834 6944 3836
rect 6648 3782 6694 3834
rect 6694 3782 6704 3834
rect 6728 3782 6758 3834
rect 6758 3782 6770 3834
rect 6770 3782 6784 3834
rect 6808 3782 6822 3834
rect 6822 3782 6834 3834
rect 6834 3782 6864 3834
rect 6888 3782 6898 3834
rect 6898 3782 6944 3834
rect 6648 3780 6704 3782
rect 6728 3780 6784 3782
rect 6808 3780 6864 3782
rect 6888 3780 6944 3782
rect 9678 5228 9734 5264
rect 9678 5208 9680 5228
rect 9680 5208 9732 5228
rect 9732 5208 9734 5228
rect 7308 3290 7364 3292
rect 7388 3290 7444 3292
rect 7468 3290 7524 3292
rect 7548 3290 7604 3292
rect 7308 3238 7354 3290
rect 7354 3238 7364 3290
rect 7388 3238 7418 3290
rect 7418 3238 7430 3290
rect 7430 3238 7444 3290
rect 7468 3238 7482 3290
rect 7482 3238 7494 3290
rect 7494 3238 7524 3290
rect 7548 3238 7558 3290
rect 7558 3238 7604 3290
rect 7308 3236 7364 3238
rect 7388 3236 7444 3238
rect 7468 3236 7524 3238
rect 7548 3236 7604 3238
rect 10506 9580 10562 9616
rect 14898 15258 14954 15260
rect 14978 15258 15034 15260
rect 15058 15258 15114 15260
rect 15138 15258 15194 15260
rect 14898 15206 14944 15258
rect 14944 15206 14954 15258
rect 14978 15206 15008 15258
rect 15008 15206 15020 15258
rect 15020 15206 15034 15258
rect 15058 15206 15072 15258
rect 15072 15206 15084 15258
rect 15084 15206 15114 15258
rect 15138 15206 15148 15258
rect 15148 15206 15194 15258
rect 14898 15204 14954 15206
rect 14978 15204 15034 15206
rect 15058 15204 15114 15206
rect 15138 15204 15194 15206
rect 14238 14714 14294 14716
rect 14318 14714 14374 14716
rect 14398 14714 14454 14716
rect 14478 14714 14534 14716
rect 14238 14662 14284 14714
rect 14284 14662 14294 14714
rect 14318 14662 14348 14714
rect 14348 14662 14360 14714
rect 14360 14662 14374 14714
rect 14398 14662 14412 14714
rect 14412 14662 14424 14714
rect 14424 14662 14454 14714
rect 14478 14662 14488 14714
rect 14488 14662 14534 14714
rect 14238 14660 14294 14662
rect 14318 14660 14374 14662
rect 14398 14660 14454 14662
rect 14478 14660 14534 14662
rect 14898 14170 14954 14172
rect 14978 14170 15034 14172
rect 15058 14170 15114 14172
rect 15138 14170 15194 14172
rect 14898 14118 14944 14170
rect 14944 14118 14954 14170
rect 14978 14118 15008 14170
rect 15008 14118 15020 14170
rect 15020 14118 15034 14170
rect 15058 14118 15072 14170
rect 15072 14118 15084 14170
rect 15084 14118 15114 14170
rect 15138 14118 15148 14170
rect 15148 14118 15194 14170
rect 14898 14116 14954 14118
rect 14978 14116 15034 14118
rect 15058 14116 15114 14118
rect 15138 14116 15194 14118
rect 14238 13626 14294 13628
rect 14318 13626 14374 13628
rect 14398 13626 14454 13628
rect 14478 13626 14534 13628
rect 14238 13574 14284 13626
rect 14284 13574 14294 13626
rect 14318 13574 14348 13626
rect 14348 13574 14360 13626
rect 14360 13574 14374 13626
rect 14398 13574 14412 13626
rect 14412 13574 14424 13626
rect 14424 13574 14454 13626
rect 14478 13574 14488 13626
rect 14488 13574 14534 13626
rect 14238 13572 14294 13574
rect 14318 13572 14374 13574
rect 14398 13572 14454 13574
rect 14478 13572 14534 13574
rect 14898 13082 14954 13084
rect 14978 13082 15034 13084
rect 15058 13082 15114 13084
rect 15138 13082 15194 13084
rect 14898 13030 14944 13082
rect 14944 13030 14954 13082
rect 14978 13030 15008 13082
rect 15008 13030 15020 13082
rect 15020 13030 15034 13082
rect 15058 13030 15072 13082
rect 15072 13030 15084 13082
rect 15084 13030 15114 13082
rect 15138 13030 15148 13082
rect 15148 13030 15194 13082
rect 14898 13028 14954 13030
rect 14978 13028 15034 13030
rect 15058 13028 15114 13030
rect 15138 13028 15194 13030
rect 14238 12538 14294 12540
rect 14318 12538 14374 12540
rect 14398 12538 14454 12540
rect 14478 12538 14534 12540
rect 14238 12486 14284 12538
rect 14284 12486 14294 12538
rect 14318 12486 14348 12538
rect 14348 12486 14360 12538
rect 14360 12486 14374 12538
rect 14398 12486 14412 12538
rect 14412 12486 14424 12538
rect 14424 12486 14454 12538
rect 14478 12486 14488 12538
rect 14488 12486 14534 12538
rect 14238 12484 14294 12486
rect 14318 12484 14374 12486
rect 14398 12484 14454 12486
rect 14478 12484 14534 12486
rect 14238 11450 14294 11452
rect 14318 11450 14374 11452
rect 14398 11450 14454 11452
rect 14478 11450 14534 11452
rect 14238 11398 14284 11450
rect 14284 11398 14294 11450
rect 14318 11398 14348 11450
rect 14348 11398 14360 11450
rect 14360 11398 14374 11450
rect 14398 11398 14412 11450
rect 14412 11398 14424 11450
rect 14424 11398 14454 11450
rect 14478 11398 14488 11450
rect 14488 11398 14534 11450
rect 14238 11396 14294 11398
rect 14318 11396 14374 11398
rect 14398 11396 14454 11398
rect 14478 11396 14534 11398
rect 14898 11994 14954 11996
rect 14978 11994 15034 11996
rect 15058 11994 15114 11996
rect 15138 11994 15194 11996
rect 14898 11942 14944 11994
rect 14944 11942 14954 11994
rect 14978 11942 15008 11994
rect 15008 11942 15020 11994
rect 15020 11942 15034 11994
rect 15058 11942 15072 11994
rect 15072 11942 15084 11994
rect 15084 11942 15114 11994
rect 15138 11942 15148 11994
rect 15148 11942 15194 11994
rect 14898 11940 14954 11942
rect 14978 11940 15034 11942
rect 15058 11940 15114 11942
rect 15138 11940 15194 11942
rect 10506 9560 10508 9580
rect 10508 9560 10560 9580
rect 10560 9560 10562 9580
rect 10443 9274 10499 9276
rect 10523 9274 10579 9276
rect 10603 9274 10659 9276
rect 10683 9274 10739 9276
rect 10443 9222 10489 9274
rect 10489 9222 10499 9274
rect 10523 9222 10553 9274
rect 10553 9222 10565 9274
rect 10565 9222 10579 9274
rect 10603 9222 10617 9274
rect 10617 9222 10629 9274
rect 10629 9222 10659 9274
rect 10683 9222 10693 9274
rect 10693 9222 10739 9274
rect 10443 9220 10499 9222
rect 10523 9220 10579 9222
rect 10603 9220 10659 9222
rect 10683 9220 10739 9222
rect 10443 8186 10499 8188
rect 10523 8186 10579 8188
rect 10603 8186 10659 8188
rect 10683 8186 10739 8188
rect 10443 8134 10489 8186
rect 10489 8134 10499 8186
rect 10523 8134 10553 8186
rect 10553 8134 10565 8186
rect 10565 8134 10579 8186
rect 10603 8134 10617 8186
rect 10617 8134 10629 8186
rect 10629 8134 10659 8186
rect 10683 8134 10693 8186
rect 10693 8134 10739 8186
rect 10443 8132 10499 8134
rect 10523 8132 10579 8134
rect 10603 8132 10659 8134
rect 10683 8132 10739 8134
rect 10443 7098 10499 7100
rect 10523 7098 10579 7100
rect 10603 7098 10659 7100
rect 10683 7098 10739 7100
rect 10443 7046 10489 7098
rect 10489 7046 10499 7098
rect 10523 7046 10553 7098
rect 10553 7046 10565 7098
rect 10565 7046 10579 7098
rect 10603 7046 10617 7098
rect 10617 7046 10629 7098
rect 10629 7046 10659 7098
rect 10683 7046 10693 7098
rect 10693 7046 10739 7098
rect 10443 7044 10499 7046
rect 10523 7044 10579 7046
rect 10603 7044 10659 7046
rect 10683 7044 10739 7046
rect 10443 6010 10499 6012
rect 10523 6010 10579 6012
rect 10603 6010 10659 6012
rect 10683 6010 10739 6012
rect 10443 5958 10489 6010
rect 10489 5958 10499 6010
rect 10523 5958 10553 6010
rect 10553 5958 10565 6010
rect 10565 5958 10579 6010
rect 10603 5958 10617 6010
rect 10617 5958 10629 6010
rect 10629 5958 10659 6010
rect 10683 5958 10693 6010
rect 10693 5958 10739 6010
rect 10443 5956 10499 5958
rect 10523 5956 10579 5958
rect 10603 5956 10659 5958
rect 10683 5956 10739 5958
rect 14238 10362 14294 10364
rect 14318 10362 14374 10364
rect 14398 10362 14454 10364
rect 14478 10362 14534 10364
rect 14238 10310 14284 10362
rect 14284 10310 14294 10362
rect 14318 10310 14348 10362
rect 14348 10310 14360 10362
rect 14360 10310 14374 10362
rect 14398 10310 14412 10362
rect 14412 10310 14424 10362
rect 14424 10310 14454 10362
rect 14478 10310 14488 10362
rect 14488 10310 14534 10362
rect 14238 10308 14294 10310
rect 14318 10308 14374 10310
rect 14398 10308 14454 10310
rect 14478 10308 14534 10310
rect 11103 8730 11159 8732
rect 11183 8730 11239 8732
rect 11263 8730 11319 8732
rect 11343 8730 11399 8732
rect 11103 8678 11149 8730
rect 11149 8678 11159 8730
rect 11183 8678 11213 8730
rect 11213 8678 11225 8730
rect 11225 8678 11239 8730
rect 11263 8678 11277 8730
rect 11277 8678 11289 8730
rect 11289 8678 11319 8730
rect 11343 8678 11353 8730
rect 11353 8678 11399 8730
rect 11103 8676 11159 8678
rect 11183 8676 11239 8678
rect 11263 8676 11319 8678
rect 11343 8676 11399 8678
rect 11103 7642 11159 7644
rect 11183 7642 11239 7644
rect 11263 7642 11319 7644
rect 11343 7642 11399 7644
rect 11103 7590 11149 7642
rect 11149 7590 11159 7642
rect 11183 7590 11213 7642
rect 11213 7590 11225 7642
rect 11225 7590 11239 7642
rect 11263 7590 11277 7642
rect 11277 7590 11289 7642
rect 11289 7590 11319 7642
rect 11343 7590 11353 7642
rect 11353 7590 11399 7642
rect 11103 7588 11159 7590
rect 11183 7588 11239 7590
rect 11263 7588 11319 7590
rect 11343 7588 11399 7590
rect 11103 6554 11159 6556
rect 11183 6554 11239 6556
rect 11263 6554 11319 6556
rect 11343 6554 11399 6556
rect 11103 6502 11149 6554
rect 11149 6502 11159 6554
rect 11183 6502 11213 6554
rect 11213 6502 11225 6554
rect 11225 6502 11239 6554
rect 11263 6502 11277 6554
rect 11277 6502 11289 6554
rect 11289 6502 11319 6554
rect 11343 6502 11353 6554
rect 11353 6502 11399 6554
rect 11103 6500 11159 6502
rect 11183 6500 11239 6502
rect 11263 6500 11319 6502
rect 11343 6500 11399 6502
rect 10443 4922 10499 4924
rect 10523 4922 10579 4924
rect 10603 4922 10659 4924
rect 10683 4922 10739 4924
rect 10443 4870 10489 4922
rect 10489 4870 10499 4922
rect 10523 4870 10553 4922
rect 10553 4870 10565 4922
rect 10565 4870 10579 4922
rect 10603 4870 10617 4922
rect 10617 4870 10629 4922
rect 10629 4870 10659 4922
rect 10683 4870 10693 4922
rect 10693 4870 10739 4922
rect 10443 4868 10499 4870
rect 10523 4868 10579 4870
rect 10603 4868 10659 4870
rect 10683 4868 10739 4870
rect 10443 3834 10499 3836
rect 10523 3834 10579 3836
rect 10603 3834 10659 3836
rect 10683 3834 10739 3836
rect 10443 3782 10489 3834
rect 10489 3782 10499 3834
rect 10523 3782 10553 3834
rect 10553 3782 10565 3834
rect 10565 3782 10579 3834
rect 10603 3782 10617 3834
rect 10617 3782 10629 3834
rect 10629 3782 10659 3834
rect 10683 3782 10693 3834
rect 10693 3782 10739 3834
rect 10443 3780 10499 3782
rect 10523 3780 10579 3782
rect 10603 3780 10659 3782
rect 10683 3780 10739 3782
rect 14238 9274 14294 9276
rect 14318 9274 14374 9276
rect 14398 9274 14454 9276
rect 14478 9274 14534 9276
rect 14238 9222 14284 9274
rect 14284 9222 14294 9274
rect 14318 9222 14348 9274
rect 14348 9222 14360 9274
rect 14360 9222 14374 9274
rect 14398 9222 14412 9274
rect 14412 9222 14424 9274
rect 14424 9222 14454 9274
rect 14478 9222 14488 9274
rect 14488 9222 14534 9274
rect 14238 9220 14294 9222
rect 14318 9220 14374 9222
rect 14398 9220 14454 9222
rect 14478 9220 14534 9222
rect 14898 10906 14954 10908
rect 14978 10906 15034 10908
rect 15058 10906 15114 10908
rect 15138 10906 15194 10908
rect 14898 10854 14944 10906
rect 14944 10854 14954 10906
rect 14978 10854 15008 10906
rect 15008 10854 15020 10906
rect 15020 10854 15034 10906
rect 15058 10854 15072 10906
rect 15072 10854 15084 10906
rect 15084 10854 15114 10906
rect 15138 10854 15148 10906
rect 15148 10854 15194 10906
rect 14898 10852 14954 10854
rect 14978 10852 15034 10854
rect 15058 10852 15114 10854
rect 15138 10852 15194 10854
rect 14898 9818 14954 9820
rect 14978 9818 15034 9820
rect 15058 9818 15114 9820
rect 15138 9818 15194 9820
rect 14898 9766 14944 9818
rect 14944 9766 14954 9818
rect 14978 9766 15008 9818
rect 15008 9766 15020 9818
rect 15020 9766 15034 9818
rect 15058 9766 15072 9818
rect 15072 9766 15084 9818
rect 15084 9766 15114 9818
rect 15138 9766 15148 9818
rect 15148 9766 15194 9818
rect 14898 9764 14954 9766
rect 14978 9764 15034 9766
rect 15058 9764 15114 9766
rect 15138 9764 15194 9766
rect 14238 8186 14294 8188
rect 14318 8186 14374 8188
rect 14398 8186 14454 8188
rect 14478 8186 14534 8188
rect 14238 8134 14284 8186
rect 14284 8134 14294 8186
rect 14318 8134 14348 8186
rect 14348 8134 14360 8186
rect 14360 8134 14374 8186
rect 14398 8134 14412 8186
rect 14412 8134 14424 8186
rect 14424 8134 14454 8186
rect 14478 8134 14488 8186
rect 14488 8134 14534 8186
rect 14238 8132 14294 8134
rect 14318 8132 14374 8134
rect 14398 8132 14454 8134
rect 14478 8132 14534 8134
rect 11103 5466 11159 5468
rect 11183 5466 11239 5468
rect 11263 5466 11319 5468
rect 11343 5466 11399 5468
rect 11103 5414 11149 5466
rect 11149 5414 11159 5466
rect 11183 5414 11213 5466
rect 11213 5414 11225 5466
rect 11225 5414 11239 5466
rect 11263 5414 11277 5466
rect 11277 5414 11289 5466
rect 11289 5414 11319 5466
rect 11343 5414 11353 5466
rect 11353 5414 11399 5466
rect 11103 5412 11159 5414
rect 11183 5412 11239 5414
rect 11263 5412 11319 5414
rect 11343 5412 11399 5414
rect 11334 5244 11336 5264
rect 11336 5244 11388 5264
rect 11388 5244 11390 5264
rect 11334 5208 11390 5244
rect 11103 4378 11159 4380
rect 11183 4378 11239 4380
rect 11263 4378 11319 4380
rect 11343 4378 11399 4380
rect 11103 4326 11149 4378
rect 11149 4326 11159 4378
rect 11183 4326 11213 4378
rect 11213 4326 11225 4378
rect 11225 4326 11239 4378
rect 11263 4326 11277 4378
rect 11277 4326 11289 4378
rect 11289 4326 11319 4378
rect 11343 4326 11353 4378
rect 11353 4326 11399 4378
rect 11103 4324 11159 4326
rect 11183 4324 11239 4326
rect 11263 4324 11319 4326
rect 11343 4324 11399 4326
rect 11103 3290 11159 3292
rect 11183 3290 11239 3292
rect 11263 3290 11319 3292
rect 11343 3290 11399 3292
rect 11103 3238 11149 3290
rect 11149 3238 11159 3290
rect 11183 3238 11213 3290
rect 11213 3238 11225 3290
rect 11225 3238 11239 3290
rect 11263 3238 11277 3290
rect 11277 3238 11289 3290
rect 11289 3238 11319 3290
rect 11343 3238 11353 3290
rect 11353 3238 11399 3290
rect 11103 3236 11159 3238
rect 11183 3236 11239 3238
rect 11263 3236 11319 3238
rect 11343 3236 11399 3238
rect 14898 8730 14954 8732
rect 14978 8730 15034 8732
rect 15058 8730 15114 8732
rect 15138 8730 15194 8732
rect 14898 8678 14944 8730
rect 14944 8678 14954 8730
rect 14978 8678 15008 8730
rect 15008 8678 15020 8730
rect 15020 8678 15034 8730
rect 15058 8678 15072 8730
rect 15072 8678 15084 8730
rect 15084 8678 15114 8730
rect 15138 8678 15148 8730
rect 15148 8678 15194 8730
rect 14898 8676 14954 8678
rect 14978 8676 15034 8678
rect 15058 8676 15114 8678
rect 15138 8676 15194 8678
rect 14898 7642 14954 7644
rect 14978 7642 15034 7644
rect 15058 7642 15114 7644
rect 15138 7642 15194 7644
rect 14898 7590 14944 7642
rect 14944 7590 14954 7642
rect 14978 7590 15008 7642
rect 15008 7590 15020 7642
rect 15020 7590 15034 7642
rect 15058 7590 15072 7642
rect 15072 7590 15084 7642
rect 15084 7590 15114 7642
rect 15138 7590 15148 7642
rect 15148 7590 15194 7642
rect 14898 7588 14954 7590
rect 14978 7588 15034 7590
rect 15058 7588 15114 7590
rect 15138 7588 15194 7590
rect 14238 7098 14294 7100
rect 14318 7098 14374 7100
rect 14398 7098 14454 7100
rect 14478 7098 14534 7100
rect 14238 7046 14284 7098
rect 14284 7046 14294 7098
rect 14318 7046 14348 7098
rect 14348 7046 14360 7098
rect 14360 7046 14374 7098
rect 14398 7046 14412 7098
rect 14412 7046 14424 7098
rect 14424 7046 14454 7098
rect 14478 7046 14488 7098
rect 14488 7046 14534 7098
rect 14238 7044 14294 7046
rect 14318 7044 14374 7046
rect 14398 7044 14454 7046
rect 14478 7044 14534 7046
rect 14238 6010 14294 6012
rect 14318 6010 14374 6012
rect 14398 6010 14454 6012
rect 14478 6010 14534 6012
rect 14238 5958 14284 6010
rect 14284 5958 14294 6010
rect 14318 5958 14348 6010
rect 14348 5958 14360 6010
rect 14360 5958 14374 6010
rect 14398 5958 14412 6010
rect 14412 5958 14424 6010
rect 14424 5958 14454 6010
rect 14478 5958 14488 6010
rect 14488 5958 14534 6010
rect 14238 5956 14294 5958
rect 14318 5956 14374 5958
rect 14398 5956 14454 5958
rect 14478 5956 14534 5958
rect 14898 6554 14954 6556
rect 14978 6554 15034 6556
rect 15058 6554 15114 6556
rect 15138 6554 15194 6556
rect 14898 6502 14944 6554
rect 14944 6502 14954 6554
rect 14978 6502 15008 6554
rect 15008 6502 15020 6554
rect 15020 6502 15034 6554
rect 15058 6502 15072 6554
rect 15072 6502 15084 6554
rect 15084 6502 15114 6554
rect 15138 6502 15148 6554
rect 15148 6502 15194 6554
rect 14898 6500 14954 6502
rect 14978 6500 15034 6502
rect 15058 6500 15114 6502
rect 15138 6500 15194 6502
rect 14898 5466 14954 5468
rect 14978 5466 15034 5468
rect 15058 5466 15114 5468
rect 15138 5466 15194 5468
rect 14898 5414 14944 5466
rect 14944 5414 14954 5466
rect 14978 5414 15008 5466
rect 15008 5414 15020 5466
rect 15020 5414 15034 5466
rect 15058 5414 15072 5466
rect 15072 5414 15084 5466
rect 15084 5414 15114 5466
rect 15138 5414 15148 5466
rect 15148 5414 15194 5466
rect 14898 5412 14954 5414
rect 14978 5412 15034 5414
rect 15058 5412 15114 5414
rect 15138 5412 15194 5414
rect 14238 4922 14294 4924
rect 14318 4922 14374 4924
rect 14398 4922 14454 4924
rect 14478 4922 14534 4924
rect 14238 4870 14284 4922
rect 14284 4870 14294 4922
rect 14318 4870 14348 4922
rect 14348 4870 14360 4922
rect 14360 4870 14374 4922
rect 14398 4870 14412 4922
rect 14412 4870 14424 4922
rect 14424 4870 14454 4922
rect 14478 4870 14488 4922
rect 14488 4870 14534 4922
rect 14238 4868 14294 4870
rect 14318 4868 14374 4870
rect 14398 4868 14454 4870
rect 14478 4868 14534 4870
rect 14898 4378 14954 4380
rect 14978 4378 15034 4380
rect 15058 4378 15114 4380
rect 15138 4378 15194 4380
rect 14898 4326 14944 4378
rect 14944 4326 14954 4378
rect 14978 4326 15008 4378
rect 15008 4326 15020 4378
rect 15020 4326 15034 4378
rect 15058 4326 15072 4378
rect 15072 4326 15084 4378
rect 15084 4326 15114 4378
rect 15138 4326 15148 4378
rect 15148 4326 15194 4378
rect 14898 4324 14954 4326
rect 14978 4324 15034 4326
rect 15058 4324 15114 4326
rect 15138 4324 15194 4326
rect 14238 3834 14294 3836
rect 14318 3834 14374 3836
rect 14398 3834 14454 3836
rect 14478 3834 14534 3836
rect 14238 3782 14284 3834
rect 14284 3782 14294 3834
rect 14318 3782 14348 3834
rect 14348 3782 14360 3834
rect 14360 3782 14374 3834
rect 14398 3782 14412 3834
rect 14412 3782 14424 3834
rect 14424 3782 14454 3834
rect 14478 3782 14488 3834
rect 14488 3782 14534 3834
rect 14238 3780 14294 3782
rect 14318 3780 14374 3782
rect 14398 3780 14454 3782
rect 14478 3780 14534 3782
rect 14898 3290 14954 3292
rect 14978 3290 15034 3292
rect 15058 3290 15114 3292
rect 15138 3290 15194 3292
rect 14898 3238 14944 3290
rect 14944 3238 14954 3290
rect 14978 3238 15008 3290
rect 15008 3238 15020 3290
rect 15020 3238 15034 3290
rect 15058 3238 15072 3290
rect 15072 3238 15084 3290
rect 15084 3238 15114 3290
rect 15138 3238 15148 3290
rect 15148 3238 15194 3290
rect 14898 3236 14954 3238
rect 14978 3236 15034 3238
rect 15058 3236 15114 3238
rect 15138 3236 15194 3238
rect 2853 2746 2909 2748
rect 2933 2746 2989 2748
rect 3013 2746 3069 2748
rect 3093 2746 3149 2748
rect 2853 2694 2899 2746
rect 2899 2694 2909 2746
rect 2933 2694 2963 2746
rect 2963 2694 2975 2746
rect 2975 2694 2989 2746
rect 3013 2694 3027 2746
rect 3027 2694 3039 2746
rect 3039 2694 3069 2746
rect 3093 2694 3103 2746
rect 3103 2694 3149 2746
rect 2853 2692 2909 2694
rect 2933 2692 2989 2694
rect 3013 2692 3069 2694
rect 3093 2692 3149 2694
rect 6648 2746 6704 2748
rect 6728 2746 6784 2748
rect 6808 2746 6864 2748
rect 6888 2746 6944 2748
rect 6648 2694 6694 2746
rect 6694 2694 6704 2746
rect 6728 2694 6758 2746
rect 6758 2694 6770 2746
rect 6770 2694 6784 2746
rect 6808 2694 6822 2746
rect 6822 2694 6834 2746
rect 6834 2694 6864 2746
rect 6888 2694 6898 2746
rect 6898 2694 6944 2746
rect 6648 2692 6704 2694
rect 6728 2692 6784 2694
rect 6808 2692 6864 2694
rect 6888 2692 6944 2694
rect 10443 2746 10499 2748
rect 10523 2746 10579 2748
rect 10603 2746 10659 2748
rect 10683 2746 10739 2748
rect 10443 2694 10489 2746
rect 10489 2694 10499 2746
rect 10523 2694 10553 2746
rect 10553 2694 10565 2746
rect 10565 2694 10579 2746
rect 10603 2694 10617 2746
rect 10617 2694 10629 2746
rect 10629 2694 10659 2746
rect 10683 2694 10693 2746
rect 10693 2694 10739 2746
rect 10443 2692 10499 2694
rect 10523 2692 10579 2694
rect 10603 2692 10659 2694
rect 10683 2692 10739 2694
rect 14238 2746 14294 2748
rect 14318 2746 14374 2748
rect 14398 2746 14454 2748
rect 14478 2746 14534 2748
rect 14238 2694 14284 2746
rect 14284 2694 14294 2746
rect 14318 2694 14348 2746
rect 14348 2694 14360 2746
rect 14360 2694 14374 2746
rect 14398 2694 14412 2746
rect 14412 2694 14424 2746
rect 14424 2694 14454 2746
rect 14478 2694 14488 2746
rect 14488 2694 14534 2746
rect 14238 2692 14294 2694
rect 14318 2692 14374 2694
rect 14398 2692 14454 2694
rect 14478 2692 14534 2694
rect 3513 2202 3569 2204
rect 3593 2202 3649 2204
rect 3673 2202 3729 2204
rect 3753 2202 3809 2204
rect 3513 2150 3559 2202
rect 3559 2150 3569 2202
rect 3593 2150 3623 2202
rect 3623 2150 3635 2202
rect 3635 2150 3649 2202
rect 3673 2150 3687 2202
rect 3687 2150 3699 2202
rect 3699 2150 3729 2202
rect 3753 2150 3763 2202
rect 3763 2150 3809 2202
rect 3513 2148 3569 2150
rect 3593 2148 3649 2150
rect 3673 2148 3729 2150
rect 3753 2148 3809 2150
rect 7308 2202 7364 2204
rect 7388 2202 7444 2204
rect 7468 2202 7524 2204
rect 7548 2202 7604 2204
rect 7308 2150 7354 2202
rect 7354 2150 7364 2202
rect 7388 2150 7418 2202
rect 7418 2150 7430 2202
rect 7430 2150 7444 2202
rect 7468 2150 7482 2202
rect 7482 2150 7494 2202
rect 7494 2150 7524 2202
rect 7548 2150 7558 2202
rect 7558 2150 7604 2202
rect 7308 2148 7364 2150
rect 7388 2148 7444 2150
rect 7468 2148 7524 2150
rect 7548 2148 7604 2150
rect 11103 2202 11159 2204
rect 11183 2202 11239 2204
rect 11263 2202 11319 2204
rect 11343 2202 11399 2204
rect 11103 2150 11149 2202
rect 11149 2150 11159 2202
rect 11183 2150 11213 2202
rect 11213 2150 11225 2202
rect 11225 2150 11239 2202
rect 11263 2150 11277 2202
rect 11277 2150 11289 2202
rect 11289 2150 11319 2202
rect 11343 2150 11353 2202
rect 11353 2150 11399 2202
rect 11103 2148 11159 2150
rect 11183 2148 11239 2150
rect 11263 2148 11319 2150
rect 11343 2148 11399 2150
rect 14898 2202 14954 2204
rect 14978 2202 15034 2204
rect 15058 2202 15114 2204
rect 15138 2202 15194 2204
rect 14898 2150 14944 2202
rect 14944 2150 14954 2202
rect 14978 2150 15008 2202
rect 15008 2150 15020 2202
rect 15020 2150 15034 2202
rect 15058 2150 15072 2202
rect 15072 2150 15084 2202
rect 15084 2150 15114 2202
rect 15138 2150 15148 2202
rect 15148 2150 15194 2202
rect 14898 2148 14954 2150
rect 14978 2148 15034 2150
rect 15058 2148 15114 2150
rect 15138 2148 15194 2150
<< metal3 >>
rect 2843 16896 3159 16897
rect 2843 16832 2849 16896
rect 2913 16832 2929 16896
rect 2993 16832 3009 16896
rect 3073 16832 3089 16896
rect 3153 16832 3159 16896
rect 2843 16831 3159 16832
rect 6638 16896 6954 16897
rect 6638 16832 6644 16896
rect 6708 16832 6724 16896
rect 6788 16832 6804 16896
rect 6868 16832 6884 16896
rect 6948 16832 6954 16896
rect 6638 16831 6954 16832
rect 10433 16896 10749 16897
rect 10433 16832 10439 16896
rect 10503 16832 10519 16896
rect 10583 16832 10599 16896
rect 10663 16832 10679 16896
rect 10743 16832 10749 16896
rect 10433 16831 10749 16832
rect 14228 16896 14544 16897
rect 14228 16832 14234 16896
rect 14298 16832 14314 16896
rect 14378 16832 14394 16896
rect 14458 16832 14474 16896
rect 14538 16832 14544 16896
rect 14228 16831 14544 16832
rect 3503 16352 3819 16353
rect 3503 16288 3509 16352
rect 3573 16288 3589 16352
rect 3653 16288 3669 16352
rect 3733 16288 3749 16352
rect 3813 16288 3819 16352
rect 3503 16287 3819 16288
rect 7298 16352 7614 16353
rect 7298 16288 7304 16352
rect 7368 16288 7384 16352
rect 7448 16288 7464 16352
rect 7528 16288 7544 16352
rect 7608 16288 7614 16352
rect 7298 16287 7614 16288
rect 11093 16352 11409 16353
rect 11093 16288 11099 16352
rect 11163 16288 11179 16352
rect 11243 16288 11259 16352
rect 11323 16288 11339 16352
rect 11403 16288 11409 16352
rect 11093 16287 11409 16288
rect 14888 16352 15204 16353
rect 14888 16288 14894 16352
rect 14958 16288 14974 16352
rect 15038 16288 15054 16352
rect 15118 16288 15134 16352
rect 15198 16288 15204 16352
rect 14888 16287 15204 16288
rect 2843 15808 3159 15809
rect 2843 15744 2849 15808
rect 2913 15744 2929 15808
rect 2993 15744 3009 15808
rect 3073 15744 3089 15808
rect 3153 15744 3159 15808
rect 2843 15743 3159 15744
rect 6638 15808 6954 15809
rect 6638 15744 6644 15808
rect 6708 15744 6724 15808
rect 6788 15744 6804 15808
rect 6868 15744 6884 15808
rect 6948 15744 6954 15808
rect 6638 15743 6954 15744
rect 10433 15808 10749 15809
rect 10433 15744 10439 15808
rect 10503 15744 10519 15808
rect 10583 15744 10599 15808
rect 10663 15744 10679 15808
rect 10743 15744 10749 15808
rect 10433 15743 10749 15744
rect 14228 15808 14544 15809
rect 14228 15744 14234 15808
rect 14298 15744 14314 15808
rect 14378 15744 14394 15808
rect 14458 15744 14474 15808
rect 14538 15744 14544 15808
rect 14228 15743 14544 15744
rect 3503 15264 3819 15265
rect 3503 15200 3509 15264
rect 3573 15200 3589 15264
rect 3653 15200 3669 15264
rect 3733 15200 3749 15264
rect 3813 15200 3819 15264
rect 3503 15199 3819 15200
rect 7298 15264 7614 15265
rect 7298 15200 7304 15264
rect 7368 15200 7384 15264
rect 7448 15200 7464 15264
rect 7528 15200 7544 15264
rect 7608 15200 7614 15264
rect 7298 15199 7614 15200
rect 11093 15264 11409 15265
rect 11093 15200 11099 15264
rect 11163 15200 11179 15264
rect 11243 15200 11259 15264
rect 11323 15200 11339 15264
rect 11403 15200 11409 15264
rect 11093 15199 11409 15200
rect 14888 15264 15204 15265
rect 14888 15200 14894 15264
rect 14958 15200 14974 15264
rect 15038 15200 15054 15264
rect 15118 15200 15134 15264
rect 15198 15200 15204 15264
rect 14888 15199 15204 15200
rect 1485 15194 1551 15197
rect 798 15192 1551 15194
rect 798 15136 1490 15192
rect 1546 15136 1551 15192
rect 798 15134 1551 15136
rect 798 15088 858 15134
rect 1485 15131 1551 15134
rect 0 14998 858 15088
rect 0 14968 800 14998
rect 2843 14720 3159 14721
rect 2843 14656 2849 14720
rect 2913 14656 2929 14720
rect 2993 14656 3009 14720
rect 3073 14656 3089 14720
rect 3153 14656 3159 14720
rect 2843 14655 3159 14656
rect 6638 14720 6954 14721
rect 6638 14656 6644 14720
rect 6708 14656 6724 14720
rect 6788 14656 6804 14720
rect 6868 14656 6884 14720
rect 6948 14656 6954 14720
rect 6638 14655 6954 14656
rect 10433 14720 10749 14721
rect 10433 14656 10439 14720
rect 10503 14656 10519 14720
rect 10583 14656 10599 14720
rect 10663 14656 10679 14720
rect 10743 14656 10749 14720
rect 10433 14655 10749 14656
rect 14228 14720 14544 14721
rect 14228 14656 14234 14720
rect 14298 14656 14314 14720
rect 14378 14656 14394 14720
rect 14458 14656 14474 14720
rect 14538 14656 14544 14720
rect 14228 14655 14544 14656
rect 3503 14176 3819 14177
rect 3503 14112 3509 14176
rect 3573 14112 3589 14176
rect 3653 14112 3669 14176
rect 3733 14112 3749 14176
rect 3813 14112 3819 14176
rect 3503 14111 3819 14112
rect 7298 14176 7614 14177
rect 7298 14112 7304 14176
rect 7368 14112 7384 14176
rect 7448 14112 7464 14176
rect 7528 14112 7544 14176
rect 7608 14112 7614 14176
rect 7298 14111 7614 14112
rect 11093 14176 11409 14177
rect 11093 14112 11099 14176
rect 11163 14112 11179 14176
rect 11243 14112 11259 14176
rect 11323 14112 11339 14176
rect 11403 14112 11409 14176
rect 11093 14111 11409 14112
rect 14888 14176 15204 14177
rect 14888 14112 14894 14176
rect 14958 14112 14974 14176
rect 15038 14112 15054 14176
rect 15118 14112 15134 14176
rect 15198 14112 15204 14176
rect 14888 14111 15204 14112
rect 2843 13632 3159 13633
rect 2843 13568 2849 13632
rect 2913 13568 2929 13632
rect 2993 13568 3009 13632
rect 3073 13568 3089 13632
rect 3153 13568 3159 13632
rect 2843 13567 3159 13568
rect 6638 13632 6954 13633
rect 6638 13568 6644 13632
rect 6708 13568 6724 13632
rect 6788 13568 6804 13632
rect 6868 13568 6884 13632
rect 6948 13568 6954 13632
rect 6638 13567 6954 13568
rect 10433 13632 10749 13633
rect 10433 13568 10439 13632
rect 10503 13568 10519 13632
rect 10583 13568 10599 13632
rect 10663 13568 10679 13632
rect 10743 13568 10749 13632
rect 10433 13567 10749 13568
rect 14228 13632 14544 13633
rect 14228 13568 14234 13632
rect 14298 13568 14314 13632
rect 14378 13568 14394 13632
rect 14458 13568 14474 13632
rect 14538 13568 14544 13632
rect 14228 13567 14544 13568
rect 3503 13088 3819 13089
rect 3503 13024 3509 13088
rect 3573 13024 3589 13088
rect 3653 13024 3669 13088
rect 3733 13024 3749 13088
rect 3813 13024 3819 13088
rect 3503 13023 3819 13024
rect 7298 13088 7614 13089
rect 7298 13024 7304 13088
rect 7368 13024 7384 13088
rect 7448 13024 7464 13088
rect 7528 13024 7544 13088
rect 7608 13024 7614 13088
rect 7298 13023 7614 13024
rect 11093 13088 11409 13089
rect 11093 13024 11099 13088
rect 11163 13024 11179 13088
rect 11243 13024 11259 13088
rect 11323 13024 11339 13088
rect 11403 13024 11409 13088
rect 11093 13023 11409 13024
rect 14888 13088 15204 13089
rect 14888 13024 14894 13088
rect 14958 13024 14974 13088
rect 15038 13024 15054 13088
rect 15118 13024 15134 13088
rect 15198 13024 15204 13088
rect 14888 13023 15204 13024
rect 2843 12544 3159 12545
rect 2843 12480 2849 12544
rect 2913 12480 2929 12544
rect 2993 12480 3009 12544
rect 3073 12480 3089 12544
rect 3153 12480 3159 12544
rect 2843 12479 3159 12480
rect 6638 12544 6954 12545
rect 6638 12480 6644 12544
rect 6708 12480 6724 12544
rect 6788 12480 6804 12544
rect 6868 12480 6884 12544
rect 6948 12480 6954 12544
rect 6638 12479 6954 12480
rect 10433 12544 10749 12545
rect 10433 12480 10439 12544
rect 10503 12480 10519 12544
rect 10583 12480 10599 12544
rect 10663 12480 10679 12544
rect 10743 12480 10749 12544
rect 10433 12479 10749 12480
rect 14228 12544 14544 12545
rect 14228 12480 14234 12544
rect 14298 12480 14314 12544
rect 14378 12480 14394 12544
rect 14458 12480 14474 12544
rect 14538 12480 14544 12544
rect 14228 12479 14544 12480
rect 3503 12000 3819 12001
rect 3503 11936 3509 12000
rect 3573 11936 3589 12000
rect 3653 11936 3669 12000
rect 3733 11936 3749 12000
rect 3813 11936 3819 12000
rect 3503 11935 3819 11936
rect 7298 12000 7614 12001
rect 7298 11936 7304 12000
rect 7368 11936 7384 12000
rect 7448 11936 7464 12000
rect 7528 11936 7544 12000
rect 7608 11936 7614 12000
rect 7298 11935 7614 11936
rect 11093 12000 11409 12001
rect 11093 11936 11099 12000
rect 11163 11936 11179 12000
rect 11243 11936 11259 12000
rect 11323 11936 11339 12000
rect 11403 11936 11409 12000
rect 11093 11935 11409 11936
rect 14888 12000 15204 12001
rect 14888 11936 14894 12000
rect 14958 11936 14974 12000
rect 15038 11936 15054 12000
rect 15118 11936 15134 12000
rect 15198 11936 15204 12000
rect 14888 11935 15204 11936
rect 13670 11596 13676 11660
rect 13740 11658 13746 11660
rect 16630 11658 17430 11688
rect 13740 11598 17430 11658
rect 13740 11596 13746 11598
rect 16630 11568 17430 11598
rect 2843 11456 3159 11457
rect 2843 11392 2849 11456
rect 2913 11392 2929 11456
rect 2993 11392 3009 11456
rect 3073 11392 3089 11456
rect 3153 11392 3159 11456
rect 2843 11391 3159 11392
rect 6638 11456 6954 11457
rect 6638 11392 6644 11456
rect 6708 11392 6724 11456
rect 6788 11392 6804 11456
rect 6868 11392 6884 11456
rect 6948 11392 6954 11456
rect 6638 11391 6954 11392
rect 10433 11456 10749 11457
rect 10433 11392 10439 11456
rect 10503 11392 10519 11456
rect 10583 11392 10599 11456
rect 10663 11392 10679 11456
rect 10743 11392 10749 11456
rect 10433 11391 10749 11392
rect 14228 11456 14544 11457
rect 14228 11392 14234 11456
rect 14298 11392 14314 11456
rect 14378 11392 14394 11456
rect 14458 11392 14474 11456
rect 14538 11392 14544 11456
rect 14228 11391 14544 11392
rect 3503 10912 3819 10913
rect 3503 10848 3509 10912
rect 3573 10848 3589 10912
rect 3653 10848 3669 10912
rect 3733 10848 3749 10912
rect 3813 10848 3819 10912
rect 3503 10847 3819 10848
rect 7298 10912 7614 10913
rect 7298 10848 7304 10912
rect 7368 10848 7384 10912
rect 7448 10848 7464 10912
rect 7528 10848 7544 10912
rect 7608 10848 7614 10912
rect 7298 10847 7614 10848
rect 11093 10912 11409 10913
rect 11093 10848 11099 10912
rect 11163 10848 11179 10912
rect 11243 10848 11259 10912
rect 11323 10848 11339 10912
rect 11403 10848 11409 10912
rect 11093 10847 11409 10848
rect 14888 10912 15204 10913
rect 14888 10848 14894 10912
rect 14958 10848 14974 10912
rect 15038 10848 15054 10912
rect 15118 10848 15134 10912
rect 15198 10848 15204 10912
rect 14888 10847 15204 10848
rect 2843 10368 3159 10369
rect 2843 10304 2849 10368
rect 2913 10304 2929 10368
rect 2993 10304 3009 10368
rect 3073 10304 3089 10368
rect 3153 10304 3159 10368
rect 2843 10303 3159 10304
rect 6638 10368 6954 10369
rect 6638 10304 6644 10368
rect 6708 10304 6724 10368
rect 6788 10304 6804 10368
rect 6868 10304 6884 10368
rect 6948 10304 6954 10368
rect 6638 10303 6954 10304
rect 10433 10368 10749 10369
rect 10433 10304 10439 10368
rect 10503 10304 10519 10368
rect 10583 10304 10599 10368
rect 10663 10304 10679 10368
rect 10743 10304 10749 10368
rect 10433 10303 10749 10304
rect 14228 10368 14544 10369
rect 14228 10304 14234 10368
rect 14298 10304 14314 10368
rect 14378 10304 14394 10368
rect 14458 10304 14474 10368
rect 14538 10304 14544 10368
rect 14228 10303 14544 10304
rect 3503 9824 3819 9825
rect 3503 9760 3509 9824
rect 3573 9760 3589 9824
rect 3653 9760 3669 9824
rect 3733 9760 3749 9824
rect 3813 9760 3819 9824
rect 3503 9759 3819 9760
rect 7298 9824 7614 9825
rect 7298 9760 7304 9824
rect 7368 9760 7384 9824
rect 7448 9760 7464 9824
rect 7528 9760 7544 9824
rect 7608 9760 7614 9824
rect 7298 9759 7614 9760
rect 11093 9824 11409 9825
rect 11093 9760 11099 9824
rect 11163 9760 11179 9824
rect 11243 9760 11259 9824
rect 11323 9760 11339 9824
rect 11403 9760 11409 9824
rect 11093 9759 11409 9760
rect 14888 9824 15204 9825
rect 14888 9760 14894 9824
rect 14958 9760 14974 9824
rect 15038 9760 15054 9824
rect 15118 9760 15134 9824
rect 15198 9760 15204 9824
rect 14888 9759 15204 9760
rect 10501 9618 10567 9621
rect 13670 9618 13676 9620
rect 10501 9616 13676 9618
rect 10501 9560 10506 9616
rect 10562 9560 13676 9616
rect 10501 9558 13676 9560
rect 10501 9555 10567 9558
rect 13670 9556 13676 9558
rect 13740 9556 13746 9620
rect 2843 9280 3159 9281
rect 2843 9216 2849 9280
rect 2913 9216 2929 9280
rect 2993 9216 3009 9280
rect 3073 9216 3089 9280
rect 3153 9216 3159 9280
rect 2843 9215 3159 9216
rect 6638 9280 6954 9281
rect 6638 9216 6644 9280
rect 6708 9216 6724 9280
rect 6788 9216 6804 9280
rect 6868 9216 6884 9280
rect 6948 9216 6954 9280
rect 6638 9215 6954 9216
rect 10433 9280 10749 9281
rect 10433 9216 10439 9280
rect 10503 9216 10519 9280
rect 10583 9216 10599 9280
rect 10663 9216 10679 9280
rect 10743 9216 10749 9280
rect 10433 9215 10749 9216
rect 14228 9280 14544 9281
rect 14228 9216 14234 9280
rect 14298 9216 14314 9280
rect 14378 9216 14394 9280
rect 14458 9216 14474 9280
rect 14538 9216 14544 9280
rect 14228 9215 14544 9216
rect 5441 9074 5507 9077
rect 9581 9074 9647 9077
rect 5441 9072 9647 9074
rect 5441 9016 5446 9072
rect 5502 9016 9586 9072
rect 9642 9016 9647 9072
rect 5441 9014 9647 9016
rect 5441 9011 5507 9014
rect 9581 9011 9647 9014
rect 3503 8736 3819 8737
rect 3503 8672 3509 8736
rect 3573 8672 3589 8736
rect 3653 8672 3669 8736
rect 3733 8672 3749 8736
rect 3813 8672 3819 8736
rect 3503 8671 3819 8672
rect 7298 8736 7614 8737
rect 7298 8672 7304 8736
rect 7368 8672 7384 8736
rect 7448 8672 7464 8736
rect 7528 8672 7544 8736
rect 7608 8672 7614 8736
rect 7298 8671 7614 8672
rect 11093 8736 11409 8737
rect 11093 8672 11099 8736
rect 11163 8672 11179 8736
rect 11243 8672 11259 8736
rect 11323 8672 11339 8736
rect 11403 8672 11409 8736
rect 11093 8671 11409 8672
rect 14888 8736 15204 8737
rect 14888 8672 14894 8736
rect 14958 8672 14974 8736
rect 15038 8672 15054 8736
rect 15118 8672 15134 8736
rect 15198 8672 15204 8736
rect 14888 8671 15204 8672
rect 2843 8192 3159 8193
rect 2843 8128 2849 8192
rect 2913 8128 2929 8192
rect 2993 8128 3009 8192
rect 3073 8128 3089 8192
rect 3153 8128 3159 8192
rect 2843 8127 3159 8128
rect 6638 8192 6954 8193
rect 6638 8128 6644 8192
rect 6708 8128 6724 8192
rect 6788 8128 6804 8192
rect 6868 8128 6884 8192
rect 6948 8128 6954 8192
rect 6638 8127 6954 8128
rect 10433 8192 10749 8193
rect 10433 8128 10439 8192
rect 10503 8128 10519 8192
rect 10583 8128 10599 8192
rect 10663 8128 10679 8192
rect 10743 8128 10749 8192
rect 10433 8127 10749 8128
rect 14228 8192 14544 8193
rect 14228 8128 14234 8192
rect 14298 8128 14314 8192
rect 14378 8128 14394 8192
rect 14458 8128 14474 8192
rect 14538 8128 14544 8192
rect 14228 8127 14544 8128
rect 3503 7648 3819 7649
rect 3503 7584 3509 7648
rect 3573 7584 3589 7648
rect 3653 7584 3669 7648
rect 3733 7584 3749 7648
rect 3813 7584 3819 7648
rect 3503 7583 3819 7584
rect 7298 7648 7614 7649
rect 7298 7584 7304 7648
rect 7368 7584 7384 7648
rect 7448 7584 7464 7648
rect 7528 7584 7544 7648
rect 7608 7584 7614 7648
rect 7298 7583 7614 7584
rect 11093 7648 11409 7649
rect 11093 7584 11099 7648
rect 11163 7584 11179 7648
rect 11243 7584 11259 7648
rect 11323 7584 11339 7648
rect 11403 7584 11409 7648
rect 11093 7583 11409 7584
rect 14888 7648 15204 7649
rect 14888 7584 14894 7648
rect 14958 7584 14974 7648
rect 15038 7584 15054 7648
rect 15118 7584 15134 7648
rect 15198 7584 15204 7648
rect 14888 7583 15204 7584
rect 2843 7104 3159 7105
rect 2843 7040 2849 7104
rect 2913 7040 2929 7104
rect 2993 7040 3009 7104
rect 3073 7040 3089 7104
rect 3153 7040 3159 7104
rect 2843 7039 3159 7040
rect 6638 7104 6954 7105
rect 6638 7040 6644 7104
rect 6708 7040 6724 7104
rect 6788 7040 6804 7104
rect 6868 7040 6884 7104
rect 6948 7040 6954 7104
rect 6638 7039 6954 7040
rect 10433 7104 10749 7105
rect 10433 7040 10439 7104
rect 10503 7040 10519 7104
rect 10583 7040 10599 7104
rect 10663 7040 10679 7104
rect 10743 7040 10749 7104
rect 10433 7039 10749 7040
rect 14228 7104 14544 7105
rect 14228 7040 14234 7104
rect 14298 7040 14314 7104
rect 14378 7040 14394 7104
rect 14458 7040 14474 7104
rect 14538 7040 14544 7104
rect 14228 7039 14544 7040
rect 3503 6560 3819 6561
rect 3503 6496 3509 6560
rect 3573 6496 3589 6560
rect 3653 6496 3669 6560
rect 3733 6496 3749 6560
rect 3813 6496 3819 6560
rect 3503 6495 3819 6496
rect 7298 6560 7614 6561
rect 7298 6496 7304 6560
rect 7368 6496 7384 6560
rect 7448 6496 7464 6560
rect 7528 6496 7544 6560
rect 7608 6496 7614 6560
rect 7298 6495 7614 6496
rect 11093 6560 11409 6561
rect 11093 6496 11099 6560
rect 11163 6496 11179 6560
rect 11243 6496 11259 6560
rect 11323 6496 11339 6560
rect 11403 6496 11409 6560
rect 11093 6495 11409 6496
rect 14888 6560 15204 6561
rect 14888 6496 14894 6560
rect 14958 6496 14974 6560
rect 15038 6496 15054 6560
rect 15118 6496 15134 6560
rect 15198 6496 15204 6560
rect 14888 6495 15204 6496
rect 2843 6016 3159 6017
rect 2843 5952 2849 6016
rect 2913 5952 2929 6016
rect 2993 5952 3009 6016
rect 3073 5952 3089 6016
rect 3153 5952 3159 6016
rect 2843 5951 3159 5952
rect 6638 6016 6954 6017
rect 6638 5952 6644 6016
rect 6708 5952 6724 6016
rect 6788 5952 6804 6016
rect 6868 5952 6884 6016
rect 6948 5952 6954 6016
rect 6638 5951 6954 5952
rect 10433 6016 10749 6017
rect 10433 5952 10439 6016
rect 10503 5952 10519 6016
rect 10583 5952 10599 6016
rect 10663 5952 10679 6016
rect 10743 5952 10749 6016
rect 10433 5951 10749 5952
rect 14228 6016 14544 6017
rect 14228 5952 14234 6016
rect 14298 5952 14314 6016
rect 14378 5952 14394 6016
rect 14458 5952 14474 6016
rect 14538 5952 14544 6016
rect 14228 5951 14544 5952
rect 3503 5472 3819 5473
rect 3503 5408 3509 5472
rect 3573 5408 3589 5472
rect 3653 5408 3669 5472
rect 3733 5408 3749 5472
rect 3813 5408 3819 5472
rect 3503 5407 3819 5408
rect 7298 5472 7614 5473
rect 7298 5408 7304 5472
rect 7368 5408 7384 5472
rect 7448 5408 7464 5472
rect 7528 5408 7544 5472
rect 7608 5408 7614 5472
rect 7298 5407 7614 5408
rect 11093 5472 11409 5473
rect 11093 5408 11099 5472
rect 11163 5408 11179 5472
rect 11243 5408 11259 5472
rect 11323 5408 11339 5472
rect 11403 5408 11409 5472
rect 11093 5407 11409 5408
rect 14888 5472 15204 5473
rect 14888 5408 14894 5472
rect 14958 5408 14974 5472
rect 15038 5408 15054 5472
rect 15118 5408 15134 5472
rect 15198 5408 15204 5472
rect 14888 5407 15204 5408
rect 9673 5266 9739 5269
rect 11329 5266 11395 5269
rect 9673 5264 11395 5266
rect 9673 5208 9678 5264
rect 9734 5208 11334 5264
rect 11390 5208 11395 5264
rect 9673 5206 11395 5208
rect 9673 5203 9739 5206
rect 11329 5203 11395 5206
rect 2843 4928 3159 4929
rect 2843 4864 2849 4928
rect 2913 4864 2929 4928
rect 2993 4864 3009 4928
rect 3073 4864 3089 4928
rect 3153 4864 3159 4928
rect 2843 4863 3159 4864
rect 6638 4928 6954 4929
rect 6638 4864 6644 4928
rect 6708 4864 6724 4928
rect 6788 4864 6804 4928
rect 6868 4864 6884 4928
rect 6948 4864 6954 4928
rect 6638 4863 6954 4864
rect 10433 4928 10749 4929
rect 10433 4864 10439 4928
rect 10503 4864 10519 4928
rect 10583 4864 10599 4928
rect 10663 4864 10679 4928
rect 10743 4864 10749 4928
rect 10433 4863 10749 4864
rect 14228 4928 14544 4929
rect 14228 4864 14234 4928
rect 14298 4864 14314 4928
rect 14378 4864 14394 4928
rect 14458 4864 14474 4928
rect 14538 4864 14544 4928
rect 14228 4863 14544 4864
rect 3503 4384 3819 4385
rect 3503 4320 3509 4384
rect 3573 4320 3589 4384
rect 3653 4320 3669 4384
rect 3733 4320 3749 4384
rect 3813 4320 3819 4384
rect 3503 4319 3819 4320
rect 7298 4384 7614 4385
rect 7298 4320 7304 4384
rect 7368 4320 7384 4384
rect 7448 4320 7464 4384
rect 7528 4320 7544 4384
rect 7608 4320 7614 4384
rect 7298 4319 7614 4320
rect 11093 4384 11409 4385
rect 11093 4320 11099 4384
rect 11163 4320 11179 4384
rect 11243 4320 11259 4384
rect 11323 4320 11339 4384
rect 11403 4320 11409 4384
rect 11093 4319 11409 4320
rect 14888 4384 15204 4385
rect 14888 4320 14894 4384
rect 14958 4320 14974 4384
rect 15038 4320 15054 4384
rect 15118 4320 15134 4384
rect 15198 4320 15204 4384
rect 14888 4319 15204 4320
rect 2843 3840 3159 3841
rect 2843 3776 2849 3840
rect 2913 3776 2929 3840
rect 2993 3776 3009 3840
rect 3073 3776 3089 3840
rect 3153 3776 3159 3840
rect 2843 3775 3159 3776
rect 6638 3840 6954 3841
rect 6638 3776 6644 3840
rect 6708 3776 6724 3840
rect 6788 3776 6804 3840
rect 6868 3776 6884 3840
rect 6948 3776 6954 3840
rect 6638 3775 6954 3776
rect 10433 3840 10749 3841
rect 10433 3776 10439 3840
rect 10503 3776 10519 3840
rect 10583 3776 10599 3840
rect 10663 3776 10679 3840
rect 10743 3776 10749 3840
rect 10433 3775 10749 3776
rect 14228 3840 14544 3841
rect 14228 3776 14234 3840
rect 14298 3776 14314 3840
rect 14378 3776 14394 3840
rect 14458 3776 14474 3840
rect 14538 3776 14544 3840
rect 14228 3775 14544 3776
rect 3503 3296 3819 3297
rect 3503 3232 3509 3296
rect 3573 3232 3589 3296
rect 3653 3232 3669 3296
rect 3733 3232 3749 3296
rect 3813 3232 3819 3296
rect 3503 3231 3819 3232
rect 7298 3296 7614 3297
rect 7298 3232 7304 3296
rect 7368 3232 7384 3296
rect 7448 3232 7464 3296
rect 7528 3232 7544 3296
rect 7608 3232 7614 3296
rect 7298 3231 7614 3232
rect 11093 3296 11409 3297
rect 11093 3232 11099 3296
rect 11163 3232 11179 3296
rect 11243 3232 11259 3296
rect 11323 3232 11339 3296
rect 11403 3232 11409 3296
rect 11093 3231 11409 3232
rect 14888 3296 15204 3297
rect 14888 3232 14894 3296
rect 14958 3232 14974 3296
rect 15038 3232 15054 3296
rect 15118 3232 15134 3296
rect 15198 3232 15204 3296
rect 14888 3231 15204 3232
rect 2843 2752 3159 2753
rect 2843 2688 2849 2752
rect 2913 2688 2929 2752
rect 2993 2688 3009 2752
rect 3073 2688 3089 2752
rect 3153 2688 3159 2752
rect 2843 2687 3159 2688
rect 6638 2752 6954 2753
rect 6638 2688 6644 2752
rect 6708 2688 6724 2752
rect 6788 2688 6804 2752
rect 6868 2688 6884 2752
rect 6948 2688 6954 2752
rect 6638 2687 6954 2688
rect 10433 2752 10749 2753
rect 10433 2688 10439 2752
rect 10503 2688 10519 2752
rect 10583 2688 10599 2752
rect 10663 2688 10679 2752
rect 10743 2688 10749 2752
rect 10433 2687 10749 2688
rect 14228 2752 14544 2753
rect 14228 2688 14234 2752
rect 14298 2688 14314 2752
rect 14378 2688 14394 2752
rect 14458 2688 14474 2752
rect 14538 2688 14544 2752
rect 14228 2687 14544 2688
rect 3503 2208 3819 2209
rect 3503 2144 3509 2208
rect 3573 2144 3589 2208
rect 3653 2144 3669 2208
rect 3733 2144 3749 2208
rect 3813 2144 3819 2208
rect 3503 2143 3819 2144
rect 7298 2208 7614 2209
rect 7298 2144 7304 2208
rect 7368 2144 7384 2208
rect 7448 2144 7464 2208
rect 7528 2144 7544 2208
rect 7608 2144 7614 2208
rect 7298 2143 7614 2144
rect 11093 2208 11409 2209
rect 11093 2144 11099 2208
rect 11163 2144 11179 2208
rect 11243 2144 11259 2208
rect 11323 2144 11339 2208
rect 11403 2144 11409 2208
rect 11093 2143 11409 2144
rect 14888 2208 15204 2209
rect 14888 2144 14894 2208
rect 14958 2144 14974 2208
rect 15038 2144 15054 2208
rect 15118 2144 15134 2208
rect 15198 2144 15204 2208
rect 14888 2143 15204 2144
<< via3 >>
rect 2849 16892 2913 16896
rect 2849 16836 2853 16892
rect 2853 16836 2909 16892
rect 2909 16836 2913 16892
rect 2849 16832 2913 16836
rect 2929 16892 2993 16896
rect 2929 16836 2933 16892
rect 2933 16836 2989 16892
rect 2989 16836 2993 16892
rect 2929 16832 2993 16836
rect 3009 16892 3073 16896
rect 3009 16836 3013 16892
rect 3013 16836 3069 16892
rect 3069 16836 3073 16892
rect 3009 16832 3073 16836
rect 3089 16892 3153 16896
rect 3089 16836 3093 16892
rect 3093 16836 3149 16892
rect 3149 16836 3153 16892
rect 3089 16832 3153 16836
rect 6644 16892 6708 16896
rect 6644 16836 6648 16892
rect 6648 16836 6704 16892
rect 6704 16836 6708 16892
rect 6644 16832 6708 16836
rect 6724 16892 6788 16896
rect 6724 16836 6728 16892
rect 6728 16836 6784 16892
rect 6784 16836 6788 16892
rect 6724 16832 6788 16836
rect 6804 16892 6868 16896
rect 6804 16836 6808 16892
rect 6808 16836 6864 16892
rect 6864 16836 6868 16892
rect 6804 16832 6868 16836
rect 6884 16892 6948 16896
rect 6884 16836 6888 16892
rect 6888 16836 6944 16892
rect 6944 16836 6948 16892
rect 6884 16832 6948 16836
rect 10439 16892 10503 16896
rect 10439 16836 10443 16892
rect 10443 16836 10499 16892
rect 10499 16836 10503 16892
rect 10439 16832 10503 16836
rect 10519 16892 10583 16896
rect 10519 16836 10523 16892
rect 10523 16836 10579 16892
rect 10579 16836 10583 16892
rect 10519 16832 10583 16836
rect 10599 16892 10663 16896
rect 10599 16836 10603 16892
rect 10603 16836 10659 16892
rect 10659 16836 10663 16892
rect 10599 16832 10663 16836
rect 10679 16892 10743 16896
rect 10679 16836 10683 16892
rect 10683 16836 10739 16892
rect 10739 16836 10743 16892
rect 10679 16832 10743 16836
rect 14234 16892 14298 16896
rect 14234 16836 14238 16892
rect 14238 16836 14294 16892
rect 14294 16836 14298 16892
rect 14234 16832 14298 16836
rect 14314 16892 14378 16896
rect 14314 16836 14318 16892
rect 14318 16836 14374 16892
rect 14374 16836 14378 16892
rect 14314 16832 14378 16836
rect 14394 16892 14458 16896
rect 14394 16836 14398 16892
rect 14398 16836 14454 16892
rect 14454 16836 14458 16892
rect 14394 16832 14458 16836
rect 14474 16892 14538 16896
rect 14474 16836 14478 16892
rect 14478 16836 14534 16892
rect 14534 16836 14538 16892
rect 14474 16832 14538 16836
rect 3509 16348 3573 16352
rect 3509 16292 3513 16348
rect 3513 16292 3569 16348
rect 3569 16292 3573 16348
rect 3509 16288 3573 16292
rect 3589 16348 3653 16352
rect 3589 16292 3593 16348
rect 3593 16292 3649 16348
rect 3649 16292 3653 16348
rect 3589 16288 3653 16292
rect 3669 16348 3733 16352
rect 3669 16292 3673 16348
rect 3673 16292 3729 16348
rect 3729 16292 3733 16348
rect 3669 16288 3733 16292
rect 3749 16348 3813 16352
rect 3749 16292 3753 16348
rect 3753 16292 3809 16348
rect 3809 16292 3813 16348
rect 3749 16288 3813 16292
rect 7304 16348 7368 16352
rect 7304 16292 7308 16348
rect 7308 16292 7364 16348
rect 7364 16292 7368 16348
rect 7304 16288 7368 16292
rect 7384 16348 7448 16352
rect 7384 16292 7388 16348
rect 7388 16292 7444 16348
rect 7444 16292 7448 16348
rect 7384 16288 7448 16292
rect 7464 16348 7528 16352
rect 7464 16292 7468 16348
rect 7468 16292 7524 16348
rect 7524 16292 7528 16348
rect 7464 16288 7528 16292
rect 7544 16348 7608 16352
rect 7544 16292 7548 16348
rect 7548 16292 7604 16348
rect 7604 16292 7608 16348
rect 7544 16288 7608 16292
rect 11099 16348 11163 16352
rect 11099 16292 11103 16348
rect 11103 16292 11159 16348
rect 11159 16292 11163 16348
rect 11099 16288 11163 16292
rect 11179 16348 11243 16352
rect 11179 16292 11183 16348
rect 11183 16292 11239 16348
rect 11239 16292 11243 16348
rect 11179 16288 11243 16292
rect 11259 16348 11323 16352
rect 11259 16292 11263 16348
rect 11263 16292 11319 16348
rect 11319 16292 11323 16348
rect 11259 16288 11323 16292
rect 11339 16348 11403 16352
rect 11339 16292 11343 16348
rect 11343 16292 11399 16348
rect 11399 16292 11403 16348
rect 11339 16288 11403 16292
rect 14894 16348 14958 16352
rect 14894 16292 14898 16348
rect 14898 16292 14954 16348
rect 14954 16292 14958 16348
rect 14894 16288 14958 16292
rect 14974 16348 15038 16352
rect 14974 16292 14978 16348
rect 14978 16292 15034 16348
rect 15034 16292 15038 16348
rect 14974 16288 15038 16292
rect 15054 16348 15118 16352
rect 15054 16292 15058 16348
rect 15058 16292 15114 16348
rect 15114 16292 15118 16348
rect 15054 16288 15118 16292
rect 15134 16348 15198 16352
rect 15134 16292 15138 16348
rect 15138 16292 15194 16348
rect 15194 16292 15198 16348
rect 15134 16288 15198 16292
rect 2849 15804 2913 15808
rect 2849 15748 2853 15804
rect 2853 15748 2909 15804
rect 2909 15748 2913 15804
rect 2849 15744 2913 15748
rect 2929 15804 2993 15808
rect 2929 15748 2933 15804
rect 2933 15748 2989 15804
rect 2989 15748 2993 15804
rect 2929 15744 2993 15748
rect 3009 15804 3073 15808
rect 3009 15748 3013 15804
rect 3013 15748 3069 15804
rect 3069 15748 3073 15804
rect 3009 15744 3073 15748
rect 3089 15804 3153 15808
rect 3089 15748 3093 15804
rect 3093 15748 3149 15804
rect 3149 15748 3153 15804
rect 3089 15744 3153 15748
rect 6644 15804 6708 15808
rect 6644 15748 6648 15804
rect 6648 15748 6704 15804
rect 6704 15748 6708 15804
rect 6644 15744 6708 15748
rect 6724 15804 6788 15808
rect 6724 15748 6728 15804
rect 6728 15748 6784 15804
rect 6784 15748 6788 15804
rect 6724 15744 6788 15748
rect 6804 15804 6868 15808
rect 6804 15748 6808 15804
rect 6808 15748 6864 15804
rect 6864 15748 6868 15804
rect 6804 15744 6868 15748
rect 6884 15804 6948 15808
rect 6884 15748 6888 15804
rect 6888 15748 6944 15804
rect 6944 15748 6948 15804
rect 6884 15744 6948 15748
rect 10439 15804 10503 15808
rect 10439 15748 10443 15804
rect 10443 15748 10499 15804
rect 10499 15748 10503 15804
rect 10439 15744 10503 15748
rect 10519 15804 10583 15808
rect 10519 15748 10523 15804
rect 10523 15748 10579 15804
rect 10579 15748 10583 15804
rect 10519 15744 10583 15748
rect 10599 15804 10663 15808
rect 10599 15748 10603 15804
rect 10603 15748 10659 15804
rect 10659 15748 10663 15804
rect 10599 15744 10663 15748
rect 10679 15804 10743 15808
rect 10679 15748 10683 15804
rect 10683 15748 10739 15804
rect 10739 15748 10743 15804
rect 10679 15744 10743 15748
rect 14234 15804 14298 15808
rect 14234 15748 14238 15804
rect 14238 15748 14294 15804
rect 14294 15748 14298 15804
rect 14234 15744 14298 15748
rect 14314 15804 14378 15808
rect 14314 15748 14318 15804
rect 14318 15748 14374 15804
rect 14374 15748 14378 15804
rect 14314 15744 14378 15748
rect 14394 15804 14458 15808
rect 14394 15748 14398 15804
rect 14398 15748 14454 15804
rect 14454 15748 14458 15804
rect 14394 15744 14458 15748
rect 14474 15804 14538 15808
rect 14474 15748 14478 15804
rect 14478 15748 14534 15804
rect 14534 15748 14538 15804
rect 14474 15744 14538 15748
rect 3509 15260 3573 15264
rect 3509 15204 3513 15260
rect 3513 15204 3569 15260
rect 3569 15204 3573 15260
rect 3509 15200 3573 15204
rect 3589 15260 3653 15264
rect 3589 15204 3593 15260
rect 3593 15204 3649 15260
rect 3649 15204 3653 15260
rect 3589 15200 3653 15204
rect 3669 15260 3733 15264
rect 3669 15204 3673 15260
rect 3673 15204 3729 15260
rect 3729 15204 3733 15260
rect 3669 15200 3733 15204
rect 3749 15260 3813 15264
rect 3749 15204 3753 15260
rect 3753 15204 3809 15260
rect 3809 15204 3813 15260
rect 3749 15200 3813 15204
rect 7304 15260 7368 15264
rect 7304 15204 7308 15260
rect 7308 15204 7364 15260
rect 7364 15204 7368 15260
rect 7304 15200 7368 15204
rect 7384 15260 7448 15264
rect 7384 15204 7388 15260
rect 7388 15204 7444 15260
rect 7444 15204 7448 15260
rect 7384 15200 7448 15204
rect 7464 15260 7528 15264
rect 7464 15204 7468 15260
rect 7468 15204 7524 15260
rect 7524 15204 7528 15260
rect 7464 15200 7528 15204
rect 7544 15260 7608 15264
rect 7544 15204 7548 15260
rect 7548 15204 7604 15260
rect 7604 15204 7608 15260
rect 7544 15200 7608 15204
rect 11099 15260 11163 15264
rect 11099 15204 11103 15260
rect 11103 15204 11159 15260
rect 11159 15204 11163 15260
rect 11099 15200 11163 15204
rect 11179 15260 11243 15264
rect 11179 15204 11183 15260
rect 11183 15204 11239 15260
rect 11239 15204 11243 15260
rect 11179 15200 11243 15204
rect 11259 15260 11323 15264
rect 11259 15204 11263 15260
rect 11263 15204 11319 15260
rect 11319 15204 11323 15260
rect 11259 15200 11323 15204
rect 11339 15260 11403 15264
rect 11339 15204 11343 15260
rect 11343 15204 11399 15260
rect 11399 15204 11403 15260
rect 11339 15200 11403 15204
rect 14894 15260 14958 15264
rect 14894 15204 14898 15260
rect 14898 15204 14954 15260
rect 14954 15204 14958 15260
rect 14894 15200 14958 15204
rect 14974 15260 15038 15264
rect 14974 15204 14978 15260
rect 14978 15204 15034 15260
rect 15034 15204 15038 15260
rect 14974 15200 15038 15204
rect 15054 15260 15118 15264
rect 15054 15204 15058 15260
rect 15058 15204 15114 15260
rect 15114 15204 15118 15260
rect 15054 15200 15118 15204
rect 15134 15260 15198 15264
rect 15134 15204 15138 15260
rect 15138 15204 15194 15260
rect 15194 15204 15198 15260
rect 15134 15200 15198 15204
rect 2849 14716 2913 14720
rect 2849 14660 2853 14716
rect 2853 14660 2909 14716
rect 2909 14660 2913 14716
rect 2849 14656 2913 14660
rect 2929 14716 2993 14720
rect 2929 14660 2933 14716
rect 2933 14660 2989 14716
rect 2989 14660 2993 14716
rect 2929 14656 2993 14660
rect 3009 14716 3073 14720
rect 3009 14660 3013 14716
rect 3013 14660 3069 14716
rect 3069 14660 3073 14716
rect 3009 14656 3073 14660
rect 3089 14716 3153 14720
rect 3089 14660 3093 14716
rect 3093 14660 3149 14716
rect 3149 14660 3153 14716
rect 3089 14656 3153 14660
rect 6644 14716 6708 14720
rect 6644 14660 6648 14716
rect 6648 14660 6704 14716
rect 6704 14660 6708 14716
rect 6644 14656 6708 14660
rect 6724 14716 6788 14720
rect 6724 14660 6728 14716
rect 6728 14660 6784 14716
rect 6784 14660 6788 14716
rect 6724 14656 6788 14660
rect 6804 14716 6868 14720
rect 6804 14660 6808 14716
rect 6808 14660 6864 14716
rect 6864 14660 6868 14716
rect 6804 14656 6868 14660
rect 6884 14716 6948 14720
rect 6884 14660 6888 14716
rect 6888 14660 6944 14716
rect 6944 14660 6948 14716
rect 6884 14656 6948 14660
rect 10439 14716 10503 14720
rect 10439 14660 10443 14716
rect 10443 14660 10499 14716
rect 10499 14660 10503 14716
rect 10439 14656 10503 14660
rect 10519 14716 10583 14720
rect 10519 14660 10523 14716
rect 10523 14660 10579 14716
rect 10579 14660 10583 14716
rect 10519 14656 10583 14660
rect 10599 14716 10663 14720
rect 10599 14660 10603 14716
rect 10603 14660 10659 14716
rect 10659 14660 10663 14716
rect 10599 14656 10663 14660
rect 10679 14716 10743 14720
rect 10679 14660 10683 14716
rect 10683 14660 10739 14716
rect 10739 14660 10743 14716
rect 10679 14656 10743 14660
rect 14234 14716 14298 14720
rect 14234 14660 14238 14716
rect 14238 14660 14294 14716
rect 14294 14660 14298 14716
rect 14234 14656 14298 14660
rect 14314 14716 14378 14720
rect 14314 14660 14318 14716
rect 14318 14660 14374 14716
rect 14374 14660 14378 14716
rect 14314 14656 14378 14660
rect 14394 14716 14458 14720
rect 14394 14660 14398 14716
rect 14398 14660 14454 14716
rect 14454 14660 14458 14716
rect 14394 14656 14458 14660
rect 14474 14716 14538 14720
rect 14474 14660 14478 14716
rect 14478 14660 14534 14716
rect 14534 14660 14538 14716
rect 14474 14656 14538 14660
rect 3509 14172 3573 14176
rect 3509 14116 3513 14172
rect 3513 14116 3569 14172
rect 3569 14116 3573 14172
rect 3509 14112 3573 14116
rect 3589 14172 3653 14176
rect 3589 14116 3593 14172
rect 3593 14116 3649 14172
rect 3649 14116 3653 14172
rect 3589 14112 3653 14116
rect 3669 14172 3733 14176
rect 3669 14116 3673 14172
rect 3673 14116 3729 14172
rect 3729 14116 3733 14172
rect 3669 14112 3733 14116
rect 3749 14172 3813 14176
rect 3749 14116 3753 14172
rect 3753 14116 3809 14172
rect 3809 14116 3813 14172
rect 3749 14112 3813 14116
rect 7304 14172 7368 14176
rect 7304 14116 7308 14172
rect 7308 14116 7364 14172
rect 7364 14116 7368 14172
rect 7304 14112 7368 14116
rect 7384 14172 7448 14176
rect 7384 14116 7388 14172
rect 7388 14116 7444 14172
rect 7444 14116 7448 14172
rect 7384 14112 7448 14116
rect 7464 14172 7528 14176
rect 7464 14116 7468 14172
rect 7468 14116 7524 14172
rect 7524 14116 7528 14172
rect 7464 14112 7528 14116
rect 7544 14172 7608 14176
rect 7544 14116 7548 14172
rect 7548 14116 7604 14172
rect 7604 14116 7608 14172
rect 7544 14112 7608 14116
rect 11099 14172 11163 14176
rect 11099 14116 11103 14172
rect 11103 14116 11159 14172
rect 11159 14116 11163 14172
rect 11099 14112 11163 14116
rect 11179 14172 11243 14176
rect 11179 14116 11183 14172
rect 11183 14116 11239 14172
rect 11239 14116 11243 14172
rect 11179 14112 11243 14116
rect 11259 14172 11323 14176
rect 11259 14116 11263 14172
rect 11263 14116 11319 14172
rect 11319 14116 11323 14172
rect 11259 14112 11323 14116
rect 11339 14172 11403 14176
rect 11339 14116 11343 14172
rect 11343 14116 11399 14172
rect 11399 14116 11403 14172
rect 11339 14112 11403 14116
rect 14894 14172 14958 14176
rect 14894 14116 14898 14172
rect 14898 14116 14954 14172
rect 14954 14116 14958 14172
rect 14894 14112 14958 14116
rect 14974 14172 15038 14176
rect 14974 14116 14978 14172
rect 14978 14116 15034 14172
rect 15034 14116 15038 14172
rect 14974 14112 15038 14116
rect 15054 14172 15118 14176
rect 15054 14116 15058 14172
rect 15058 14116 15114 14172
rect 15114 14116 15118 14172
rect 15054 14112 15118 14116
rect 15134 14172 15198 14176
rect 15134 14116 15138 14172
rect 15138 14116 15194 14172
rect 15194 14116 15198 14172
rect 15134 14112 15198 14116
rect 2849 13628 2913 13632
rect 2849 13572 2853 13628
rect 2853 13572 2909 13628
rect 2909 13572 2913 13628
rect 2849 13568 2913 13572
rect 2929 13628 2993 13632
rect 2929 13572 2933 13628
rect 2933 13572 2989 13628
rect 2989 13572 2993 13628
rect 2929 13568 2993 13572
rect 3009 13628 3073 13632
rect 3009 13572 3013 13628
rect 3013 13572 3069 13628
rect 3069 13572 3073 13628
rect 3009 13568 3073 13572
rect 3089 13628 3153 13632
rect 3089 13572 3093 13628
rect 3093 13572 3149 13628
rect 3149 13572 3153 13628
rect 3089 13568 3153 13572
rect 6644 13628 6708 13632
rect 6644 13572 6648 13628
rect 6648 13572 6704 13628
rect 6704 13572 6708 13628
rect 6644 13568 6708 13572
rect 6724 13628 6788 13632
rect 6724 13572 6728 13628
rect 6728 13572 6784 13628
rect 6784 13572 6788 13628
rect 6724 13568 6788 13572
rect 6804 13628 6868 13632
rect 6804 13572 6808 13628
rect 6808 13572 6864 13628
rect 6864 13572 6868 13628
rect 6804 13568 6868 13572
rect 6884 13628 6948 13632
rect 6884 13572 6888 13628
rect 6888 13572 6944 13628
rect 6944 13572 6948 13628
rect 6884 13568 6948 13572
rect 10439 13628 10503 13632
rect 10439 13572 10443 13628
rect 10443 13572 10499 13628
rect 10499 13572 10503 13628
rect 10439 13568 10503 13572
rect 10519 13628 10583 13632
rect 10519 13572 10523 13628
rect 10523 13572 10579 13628
rect 10579 13572 10583 13628
rect 10519 13568 10583 13572
rect 10599 13628 10663 13632
rect 10599 13572 10603 13628
rect 10603 13572 10659 13628
rect 10659 13572 10663 13628
rect 10599 13568 10663 13572
rect 10679 13628 10743 13632
rect 10679 13572 10683 13628
rect 10683 13572 10739 13628
rect 10739 13572 10743 13628
rect 10679 13568 10743 13572
rect 14234 13628 14298 13632
rect 14234 13572 14238 13628
rect 14238 13572 14294 13628
rect 14294 13572 14298 13628
rect 14234 13568 14298 13572
rect 14314 13628 14378 13632
rect 14314 13572 14318 13628
rect 14318 13572 14374 13628
rect 14374 13572 14378 13628
rect 14314 13568 14378 13572
rect 14394 13628 14458 13632
rect 14394 13572 14398 13628
rect 14398 13572 14454 13628
rect 14454 13572 14458 13628
rect 14394 13568 14458 13572
rect 14474 13628 14538 13632
rect 14474 13572 14478 13628
rect 14478 13572 14534 13628
rect 14534 13572 14538 13628
rect 14474 13568 14538 13572
rect 3509 13084 3573 13088
rect 3509 13028 3513 13084
rect 3513 13028 3569 13084
rect 3569 13028 3573 13084
rect 3509 13024 3573 13028
rect 3589 13084 3653 13088
rect 3589 13028 3593 13084
rect 3593 13028 3649 13084
rect 3649 13028 3653 13084
rect 3589 13024 3653 13028
rect 3669 13084 3733 13088
rect 3669 13028 3673 13084
rect 3673 13028 3729 13084
rect 3729 13028 3733 13084
rect 3669 13024 3733 13028
rect 3749 13084 3813 13088
rect 3749 13028 3753 13084
rect 3753 13028 3809 13084
rect 3809 13028 3813 13084
rect 3749 13024 3813 13028
rect 7304 13084 7368 13088
rect 7304 13028 7308 13084
rect 7308 13028 7364 13084
rect 7364 13028 7368 13084
rect 7304 13024 7368 13028
rect 7384 13084 7448 13088
rect 7384 13028 7388 13084
rect 7388 13028 7444 13084
rect 7444 13028 7448 13084
rect 7384 13024 7448 13028
rect 7464 13084 7528 13088
rect 7464 13028 7468 13084
rect 7468 13028 7524 13084
rect 7524 13028 7528 13084
rect 7464 13024 7528 13028
rect 7544 13084 7608 13088
rect 7544 13028 7548 13084
rect 7548 13028 7604 13084
rect 7604 13028 7608 13084
rect 7544 13024 7608 13028
rect 11099 13084 11163 13088
rect 11099 13028 11103 13084
rect 11103 13028 11159 13084
rect 11159 13028 11163 13084
rect 11099 13024 11163 13028
rect 11179 13084 11243 13088
rect 11179 13028 11183 13084
rect 11183 13028 11239 13084
rect 11239 13028 11243 13084
rect 11179 13024 11243 13028
rect 11259 13084 11323 13088
rect 11259 13028 11263 13084
rect 11263 13028 11319 13084
rect 11319 13028 11323 13084
rect 11259 13024 11323 13028
rect 11339 13084 11403 13088
rect 11339 13028 11343 13084
rect 11343 13028 11399 13084
rect 11399 13028 11403 13084
rect 11339 13024 11403 13028
rect 14894 13084 14958 13088
rect 14894 13028 14898 13084
rect 14898 13028 14954 13084
rect 14954 13028 14958 13084
rect 14894 13024 14958 13028
rect 14974 13084 15038 13088
rect 14974 13028 14978 13084
rect 14978 13028 15034 13084
rect 15034 13028 15038 13084
rect 14974 13024 15038 13028
rect 15054 13084 15118 13088
rect 15054 13028 15058 13084
rect 15058 13028 15114 13084
rect 15114 13028 15118 13084
rect 15054 13024 15118 13028
rect 15134 13084 15198 13088
rect 15134 13028 15138 13084
rect 15138 13028 15194 13084
rect 15194 13028 15198 13084
rect 15134 13024 15198 13028
rect 2849 12540 2913 12544
rect 2849 12484 2853 12540
rect 2853 12484 2909 12540
rect 2909 12484 2913 12540
rect 2849 12480 2913 12484
rect 2929 12540 2993 12544
rect 2929 12484 2933 12540
rect 2933 12484 2989 12540
rect 2989 12484 2993 12540
rect 2929 12480 2993 12484
rect 3009 12540 3073 12544
rect 3009 12484 3013 12540
rect 3013 12484 3069 12540
rect 3069 12484 3073 12540
rect 3009 12480 3073 12484
rect 3089 12540 3153 12544
rect 3089 12484 3093 12540
rect 3093 12484 3149 12540
rect 3149 12484 3153 12540
rect 3089 12480 3153 12484
rect 6644 12540 6708 12544
rect 6644 12484 6648 12540
rect 6648 12484 6704 12540
rect 6704 12484 6708 12540
rect 6644 12480 6708 12484
rect 6724 12540 6788 12544
rect 6724 12484 6728 12540
rect 6728 12484 6784 12540
rect 6784 12484 6788 12540
rect 6724 12480 6788 12484
rect 6804 12540 6868 12544
rect 6804 12484 6808 12540
rect 6808 12484 6864 12540
rect 6864 12484 6868 12540
rect 6804 12480 6868 12484
rect 6884 12540 6948 12544
rect 6884 12484 6888 12540
rect 6888 12484 6944 12540
rect 6944 12484 6948 12540
rect 6884 12480 6948 12484
rect 10439 12540 10503 12544
rect 10439 12484 10443 12540
rect 10443 12484 10499 12540
rect 10499 12484 10503 12540
rect 10439 12480 10503 12484
rect 10519 12540 10583 12544
rect 10519 12484 10523 12540
rect 10523 12484 10579 12540
rect 10579 12484 10583 12540
rect 10519 12480 10583 12484
rect 10599 12540 10663 12544
rect 10599 12484 10603 12540
rect 10603 12484 10659 12540
rect 10659 12484 10663 12540
rect 10599 12480 10663 12484
rect 10679 12540 10743 12544
rect 10679 12484 10683 12540
rect 10683 12484 10739 12540
rect 10739 12484 10743 12540
rect 10679 12480 10743 12484
rect 14234 12540 14298 12544
rect 14234 12484 14238 12540
rect 14238 12484 14294 12540
rect 14294 12484 14298 12540
rect 14234 12480 14298 12484
rect 14314 12540 14378 12544
rect 14314 12484 14318 12540
rect 14318 12484 14374 12540
rect 14374 12484 14378 12540
rect 14314 12480 14378 12484
rect 14394 12540 14458 12544
rect 14394 12484 14398 12540
rect 14398 12484 14454 12540
rect 14454 12484 14458 12540
rect 14394 12480 14458 12484
rect 14474 12540 14538 12544
rect 14474 12484 14478 12540
rect 14478 12484 14534 12540
rect 14534 12484 14538 12540
rect 14474 12480 14538 12484
rect 3509 11996 3573 12000
rect 3509 11940 3513 11996
rect 3513 11940 3569 11996
rect 3569 11940 3573 11996
rect 3509 11936 3573 11940
rect 3589 11996 3653 12000
rect 3589 11940 3593 11996
rect 3593 11940 3649 11996
rect 3649 11940 3653 11996
rect 3589 11936 3653 11940
rect 3669 11996 3733 12000
rect 3669 11940 3673 11996
rect 3673 11940 3729 11996
rect 3729 11940 3733 11996
rect 3669 11936 3733 11940
rect 3749 11996 3813 12000
rect 3749 11940 3753 11996
rect 3753 11940 3809 11996
rect 3809 11940 3813 11996
rect 3749 11936 3813 11940
rect 7304 11996 7368 12000
rect 7304 11940 7308 11996
rect 7308 11940 7364 11996
rect 7364 11940 7368 11996
rect 7304 11936 7368 11940
rect 7384 11996 7448 12000
rect 7384 11940 7388 11996
rect 7388 11940 7444 11996
rect 7444 11940 7448 11996
rect 7384 11936 7448 11940
rect 7464 11996 7528 12000
rect 7464 11940 7468 11996
rect 7468 11940 7524 11996
rect 7524 11940 7528 11996
rect 7464 11936 7528 11940
rect 7544 11996 7608 12000
rect 7544 11940 7548 11996
rect 7548 11940 7604 11996
rect 7604 11940 7608 11996
rect 7544 11936 7608 11940
rect 11099 11996 11163 12000
rect 11099 11940 11103 11996
rect 11103 11940 11159 11996
rect 11159 11940 11163 11996
rect 11099 11936 11163 11940
rect 11179 11996 11243 12000
rect 11179 11940 11183 11996
rect 11183 11940 11239 11996
rect 11239 11940 11243 11996
rect 11179 11936 11243 11940
rect 11259 11996 11323 12000
rect 11259 11940 11263 11996
rect 11263 11940 11319 11996
rect 11319 11940 11323 11996
rect 11259 11936 11323 11940
rect 11339 11996 11403 12000
rect 11339 11940 11343 11996
rect 11343 11940 11399 11996
rect 11399 11940 11403 11996
rect 11339 11936 11403 11940
rect 14894 11996 14958 12000
rect 14894 11940 14898 11996
rect 14898 11940 14954 11996
rect 14954 11940 14958 11996
rect 14894 11936 14958 11940
rect 14974 11996 15038 12000
rect 14974 11940 14978 11996
rect 14978 11940 15034 11996
rect 15034 11940 15038 11996
rect 14974 11936 15038 11940
rect 15054 11996 15118 12000
rect 15054 11940 15058 11996
rect 15058 11940 15114 11996
rect 15114 11940 15118 11996
rect 15054 11936 15118 11940
rect 15134 11996 15198 12000
rect 15134 11940 15138 11996
rect 15138 11940 15194 11996
rect 15194 11940 15198 11996
rect 15134 11936 15198 11940
rect 13676 11596 13740 11660
rect 2849 11452 2913 11456
rect 2849 11396 2853 11452
rect 2853 11396 2909 11452
rect 2909 11396 2913 11452
rect 2849 11392 2913 11396
rect 2929 11452 2993 11456
rect 2929 11396 2933 11452
rect 2933 11396 2989 11452
rect 2989 11396 2993 11452
rect 2929 11392 2993 11396
rect 3009 11452 3073 11456
rect 3009 11396 3013 11452
rect 3013 11396 3069 11452
rect 3069 11396 3073 11452
rect 3009 11392 3073 11396
rect 3089 11452 3153 11456
rect 3089 11396 3093 11452
rect 3093 11396 3149 11452
rect 3149 11396 3153 11452
rect 3089 11392 3153 11396
rect 6644 11452 6708 11456
rect 6644 11396 6648 11452
rect 6648 11396 6704 11452
rect 6704 11396 6708 11452
rect 6644 11392 6708 11396
rect 6724 11452 6788 11456
rect 6724 11396 6728 11452
rect 6728 11396 6784 11452
rect 6784 11396 6788 11452
rect 6724 11392 6788 11396
rect 6804 11452 6868 11456
rect 6804 11396 6808 11452
rect 6808 11396 6864 11452
rect 6864 11396 6868 11452
rect 6804 11392 6868 11396
rect 6884 11452 6948 11456
rect 6884 11396 6888 11452
rect 6888 11396 6944 11452
rect 6944 11396 6948 11452
rect 6884 11392 6948 11396
rect 10439 11452 10503 11456
rect 10439 11396 10443 11452
rect 10443 11396 10499 11452
rect 10499 11396 10503 11452
rect 10439 11392 10503 11396
rect 10519 11452 10583 11456
rect 10519 11396 10523 11452
rect 10523 11396 10579 11452
rect 10579 11396 10583 11452
rect 10519 11392 10583 11396
rect 10599 11452 10663 11456
rect 10599 11396 10603 11452
rect 10603 11396 10659 11452
rect 10659 11396 10663 11452
rect 10599 11392 10663 11396
rect 10679 11452 10743 11456
rect 10679 11396 10683 11452
rect 10683 11396 10739 11452
rect 10739 11396 10743 11452
rect 10679 11392 10743 11396
rect 14234 11452 14298 11456
rect 14234 11396 14238 11452
rect 14238 11396 14294 11452
rect 14294 11396 14298 11452
rect 14234 11392 14298 11396
rect 14314 11452 14378 11456
rect 14314 11396 14318 11452
rect 14318 11396 14374 11452
rect 14374 11396 14378 11452
rect 14314 11392 14378 11396
rect 14394 11452 14458 11456
rect 14394 11396 14398 11452
rect 14398 11396 14454 11452
rect 14454 11396 14458 11452
rect 14394 11392 14458 11396
rect 14474 11452 14538 11456
rect 14474 11396 14478 11452
rect 14478 11396 14534 11452
rect 14534 11396 14538 11452
rect 14474 11392 14538 11396
rect 3509 10908 3573 10912
rect 3509 10852 3513 10908
rect 3513 10852 3569 10908
rect 3569 10852 3573 10908
rect 3509 10848 3573 10852
rect 3589 10908 3653 10912
rect 3589 10852 3593 10908
rect 3593 10852 3649 10908
rect 3649 10852 3653 10908
rect 3589 10848 3653 10852
rect 3669 10908 3733 10912
rect 3669 10852 3673 10908
rect 3673 10852 3729 10908
rect 3729 10852 3733 10908
rect 3669 10848 3733 10852
rect 3749 10908 3813 10912
rect 3749 10852 3753 10908
rect 3753 10852 3809 10908
rect 3809 10852 3813 10908
rect 3749 10848 3813 10852
rect 7304 10908 7368 10912
rect 7304 10852 7308 10908
rect 7308 10852 7364 10908
rect 7364 10852 7368 10908
rect 7304 10848 7368 10852
rect 7384 10908 7448 10912
rect 7384 10852 7388 10908
rect 7388 10852 7444 10908
rect 7444 10852 7448 10908
rect 7384 10848 7448 10852
rect 7464 10908 7528 10912
rect 7464 10852 7468 10908
rect 7468 10852 7524 10908
rect 7524 10852 7528 10908
rect 7464 10848 7528 10852
rect 7544 10908 7608 10912
rect 7544 10852 7548 10908
rect 7548 10852 7604 10908
rect 7604 10852 7608 10908
rect 7544 10848 7608 10852
rect 11099 10908 11163 10912
rect 11099 10852 11103 10908
rect 11103 10852 11159 10908
rect 11159 10852 11163 10908
rect 11099 10848 11163 10852
rect 11179 10908 11243 10912
rect 11179 10852 11183 10908
rect 11183 10852 11239 10908
rect 11239 10852 11243 10908
rect 11179 10848 11243 10852
rect 11259 10908 11323 10912
rect 11259 10852 11263 10908
rect 11263 10852 11319 10908
rect 11319 10852 11323 10908
rect 11259 10848 11323 10852
rect 11339 10908 11403 10912
rect 11339 10852 11343 10908
rect 11343 10852 11399 10908
rect 11399 10852 11403 10908
rect 11339 10848 11403 10852
rect 14894 10908 14958 10912
rect 14894 10852 14898 10908
rect 14898 10852 14954 10908
rect 14954 10852 14958 10908
rect 14894 10848 14958 10852
rect 14974 10908 15038 10912
rect 14974 10852 14978 10908
rect 14978 10852 15034 10908
rect 15034 10852 15038 10908
rect 14974 10848 15038 10852
rect 15054 10908 15118 10912
rect 15054 10852 15058 10908
rect 15058 10852 15114 10908
rect 15114 10852 15118 10908
rect 15054 10848 15118 10852
rect 15134 10908 15198 10912
rect 15134 10852 15138 10908
rect 15138 10852 15194 10908
rect 15194 10852 15198 10908
rect 15134 10848 15198 10852
rect 2849 10364 2913 10368
rect 2849 10308 2853 10364
rect 2853 10308 2909 10364
rect 2909 10308 2913 10364
rect 2849 10304 2913 10308
rect 2929 10364 2993 10368
rect 2929 10308 2933 10364
rect 2933 10308 2989 10364
rect 2989 10308 2993 10364
rect 2929 10304 2993 10308
rect 3009 10364 3073 10368
rect 3009 10308 3013 10364
rect 3013 10308 3069 10364
rect 3069 10308 3073 10364
rect 3009 10304 3073 10308
rect 3089 10364 3153 10368
rect 3089 10308 3093 10364
rect 3093 10308 3149 10364
rect 3149 10308 3153 10364
rect 3089 10304 3153 10308
rect 6644 10364 6708 10368
rect 6644 10308 6648 10364
rect 6648 10308 6704 10364
rect 6704 10308 6708 10364
rect 6644 10304 6708 10308
rect 6724 10364 6788 10368
rect 6724 10308 6728 10364
rect 6728 10308 6784 10364
rect 6784 10308 6788 10364
rect 6724 10304 6788 10308
rect 6804 10364 6868 10368
rect 6804 10308 6808 10364
rect 6808 10308 6864 10364
rect 6864 10308 6868 10364
rect 6804 10304 6868 10308
rect 6884 10364 6948 10368
rect 6884 10308 6888 10364
rect 6888 10308 6944 10364
rect 6944 10308 6948 10364
rect 6884 10304 6948 10308
rect 10439 10364 10503 10368
rect 10439 10308 10443 10364
rect 10443 10308 10499 10364
rect 10499 10308 10503 10364
rect 10439 10304 10503 10308
rect 10519 10364 10583 10368
rect 10519 10308 10523 10364
rect 10523 10308 10579 10364
rect 10579 10308 10583 10364
rect 10519 10304 10583 10308
rect 10599 10364 10663 10368
rect 10599 10308 10603 10364
rect 10603 10308 10659 10364
rect 10659 10308 10663 10364
rect 10599 10304 10663 10308
rect 10679 10364 10743 10368
rect 10679 10308 10683 10364
rect 10683 10308 10739 10364
rect 10739 10308 10743 10364
rect 10679 10304 10743 10308
rect 14234 10364 14298 10368
rect 14234 10308 14238 10364
rect 14238 10308 14294 10364
rect 14294 10308 14298 10364
rect 14234 10304 14298 10308
rect 14314 10364 14378 10368
rect 14314 10308 14318 10364
rect 14318 10308 14374 10364
rect 14374 10308 14378 10364
rect 14314 10304 14378 10308
rect 14394 10364 14458 10368
rect 14394 10308 14398 10364
rect 14398 10308 14454 10364
rect 14454 10308 14458 10364
rect 14394 10304 14458 10308
rect 14474 10364 14538 10368
rect 14474 10308 14478 10364
rect 14478 10308 14534 10364
rect 14534 10308 14538 10364
rect 14474 10304 14538 10308
rect 3509 9820 3573 9824
rect 3509 9764 3513 9820
rect 3513 9764 3569 9820
rect 3569 9764 3573 9820
rect 3509 9760 3573 9764
rect 3589 9820 3653 9824
rect 3589 9764 3593 9820
rect 3593 9764 3649 9820
rect 3649 9764 3653 9820
rect 3589 9760 3653 9764
rect 3669 9820 3733 9824
rect 3669 9764 3673 9820
rect 3673 9764 3729 9820
rect 3729 9764 3733 9820
rect 3669 9760 3733 9764
rect 3749 9820 3813 9824
rect 3749 9764 3753 9820
rect 3753 9764 3809 9820
rect 3809 9764 3813 9820
rect 3749 9760 3813 9764
rect 7304 9820 7368 9824
rect 7304 9764 7308 9820
rect 7308 9764 7364 9820
rect 7364 9764 7368 9820
rect 7304 9760 7368 9764
rect 7384 9820 7448 9824
rect 7384 9764 7388 9820
rect 7388 9764 7444 9820
rect 7444 9764 7448 9820
rect 7384 9760 7448 9764
rect 7464 9820 7528 9824
rect 7464 9764 7468 9820
rect 7468 9764 7524 9820
rect 7524 9764 7528 9820
rect 7464 9760 7528 9764
rect 7544 9820 7608 9824
rect 7544 9764 7548 9820
rect 7548 9764 7604 9820
rect 7604 9764 7608 9820
rect 7544 9760 7608 9764
rect 11099 9820 11163 9824
rect 11099 9764 11103 9820
rect 11103 9764 11159 9820
rect 11159 9764 11163 9820
rect 11099 9760 11163 9764
rect 11179 9820 11243 9824
rect 11179 9764 11183 9820
rect 11183 9764 11239 9820
rect 11239 9764 11243 9820
rect 11179 9760 11243 9764
rect 11259 9820 11323 9824
rect 11259 9764 11263 9820
rect 11263 9764 11319 9820
rect 11319 9764 11323 9820
rect 11259 9760 11323 9764
rect 11339 9820 11403 9824
rect 11339 9764 11343 9820
rect 11343 9764 11399 9820
rect 11399 9764 11403 9820
rect 11339 9760 11403 9764
rect 14894 9820 14958 9824
rect 14894 9764 14898 9820
rect 14898 9764 14954 9820
rect 14954 9764 14958 9820
rect 14894 9760 14958 9764
rect 14974 9820 15038 9824
rect 14974 9764 14978 9820
rect 14978 9764 15034 9820
rect 15034 9764 15038 9820
rect 14974 9760 15038 9764
rect 15054 9820 15118 9824
rect 15054 9764 15058 9820
rect 15058 9764 15114 9820
rect 15114 9764 15118 9820
rect 15054 9760 15118 9764
rect 15134 9820 15198 9824
rect 15134 9764 15138 9820
rect 15138 9764 15194 9820
rect 15194 9764 15198 9820
rect 15134 9760 15198 9764
rect 13676 9556 13740 9620
rect 2849 9276 2913 9280
rect 2849 9220 2853 9276
rect 2853 9220 2909 9276
rect 2909 9220 2913 9276
rect 2849 9216 2913 9220
rect 2929 9276 2993 9280
rect 2929 9220 2933 9276
rect 2933 9220 2989 9276
rect 2989 9220 2993 9276
rect 2929 9216 2993 9220
rect 3009 9276 3073 9280
rect 3009 9220 3013 9276
rect 3013 9220 3069 9276
rect 3069 9220 3073 9276
rect 3009 9216 3073 9220
rect 3089 9276 3153 9280
rect 3089 9220 3093 9276
rect 3093 9220 3149 9276
rect 3149 9220 3153 9276
rect 3089 9216 3153 9220
rect 6644 9276 6708 9280
rect 6644 9220 6648 9276
rect 6648 9220 6704 9276
rect 6704 9220 6708 9276
rect 6644 9216 6708 9220
rect 6724 9276 6788 9280
rect 6724 9220 6728 9276
rect 6728 9220 6784 9276
rect 6784 9220 6788 9276
rect 6724 9216 6788 9220
rect 6804 9276 6868 9280
rect 6804 9220 6808 9276
rect 6808 9220 6864 9276
rect 6864 9220 6868 9276
rect 6804 9216 6868 9220
rect 6884 9276 6948 9280
rect 6884 9220 6888 9276
rect 6888 9220 6944 9276
rect 6944 9220 6948 9276
rect 6884 9216 6948 9220
rect 10439 9276 10503 9280
rect 10439 9220 10443 9276
rect 10443 9220 10499 9276
rect 10499 9220 10503 9276
rect 10439 9216 10503 9220
rect 10519 9276 10583 9280
rect 10519 9220 10523 9276
rect 10523 9220 10579 9276
rect 10579 9220 10583 9276
rect 10519 9216 10583 9220
rect 10599 9276 10663 9280
rect 10599 9220 10603 9276
rect 10603 9220 10659 9276
rect 10659 9220 10663 9276
rect 10599 9216 10663 9220
rect 10679 9276 10743 9280
rect 10679 9220 10683 9276
rect 10683 9220 10739 9276
rect 10739 9220 10743 9276
rect 10679 9216 10743 9220
rect 14234 9276 14298 9280
rect 14234 9220 14238 9276
rect 14238 9220 14294 9276
rect 14294 9220 14298 9276
rect 14234 9216 14298 9220
rect 14314 9276 14378 9280
rect 14314 9220 14318 9276
rect 14318 9220 14374 9276
rect 14374 9220 14378 9276
rect 14314 9216 14378 9220
rect 14394 9276 14458 9280
rect 14394 9220 14398 9276
rect 14398 9220 14454 9276
rect 14454 9220 14458 9276
rect 14394 9216 14458 9220
rect 14474 9276 14538 9280
rect 14474 9220 14478 9276
rect 14478 9220 14534 9276
rect 14534 9220 14538 9276
rect 14474 9216 14538 9220
rect 3509 8732 3573 8736
rect 3509 8676 3513 8732
rect 3513 8676 3569 8732
rect 3569 8676 3573 8732
rect 3509 8672 3573 8676
rect 3589 8732 3653 8736
rect 3589 8676 3593 8732
rect 3593 8676 3649 8732
rect 3649 8676 3653 8732
rect 3589 8672 3653 8676
rect 3669 8732 3733 8736
rect 3669 8676 3673 8732
rect 3673 8676 3729 8732
rect 3729 8676 3733 8732
rect 3669 8672 3733 8676
rect 3749 8732 3813 8736
rect 3749 8676 3753 8732
rect 3753 8676 3809 8732
rect 3809 8676 3813 8732
rect 3749 8672 3813 8676
rect 7304 8732 7368 8736
rect 7304 8676 7308 8732
rect 7308 8676 7364 8732
rect 7364 8676 7368 8732
rect 7304 8672 7368 8676
rect 7384 8732 7448 8736
rect 7384 8676 7388 8732
rect 7388 8676 7444 8732
rect 7444 8676 7448 8732
rect 7384 8672 7448 8676
rect 7464 8732 7528 8736
rect 7464 8676 7468 8732
rect 7468 8676 7524 8732
rect 7524 8676 7528 8732
rect 7464 8672 7528 8676
rect 7544 8732 7608 8736
rect 7544 8676 7548 8732
rect 7548 8676 7604 8732
rect 7604 8676 7608 8732
rect 7544 8672 7608 8676
rect 11099 8732 11163 8736
rect 11099 8676 11103 8732
rect 11103 8676 11159 8732
rect 11159 8676 11163 8732
rect 11099 8672 11163 8676
rect 11179 8732 11243 8736
rect 11179 8676 11183 8732
rect 11183 8676 11239 8732
rect 11239 8676 11243 8732
rect 11179 8672 11243 8676
rect 11259 8732 11323 8736
rect 11259 8676 11263 8732
rect 11263 8676 11319 8732
rect 11319 8676 11323 8732
rect 11259 8672 11323 8676
rect 11339 8732 11403 8736
rect 11339 8676 11343 8732
rect 11343 8676 11399 8732
rect 11399 8676 11403 8732
rect 11339 8672 11403 8676
rect 14894 8732 14958 8736
rect 14894 8676 14898 8732
rect 14898 8676 14954 8732
rect 14954 8676 14958 8732
rect 14894 8672 14958 8676
rect 14974 8732 15038 8736
rect 14974 8676 14978 8732
rect 14978 8676 15034 8732
rect 15034 8676 15038 8732
rect 14974 8672 15038 8676
rect 15054 8732 15118 8736
rect 15054 8676 15058 8732
rect 15058 8676 15114 8732
rect 15114 8676 15118 8732
rect 15054 8672 15118 8676
rect 15134 8732 15198 8736
rect 15134 8676 15138 8732
rect 15138 8676 15194 8732
rect 15194 8676 15198 8732
rect 15134 8672 15198 8676
rect 2849 8188 2913 8192
rect 2849 8132 2853 8188
rect 2853 8132 2909 8188
rect 2909 8132 2913 8188
rect 2849 8128 2913 8132
rect 2929 8188 2993 8192
rect 2929 8132 2933 8188
rect 2933 8132 2989 8188
rect 2989 8132 2993 8188
rect 2929 8128 2993 8132
rect 3009 8188 3073 8192
rect 3009 8132 3013 8188
rect 3013 8132 3069 8188
rect 3069 8132 3073 8188
rect 3009 8128 3073 8132
rect 3089 8188 3153 8192
rect 3089 8132 3093 8188
rect 3093 8132 3149 8188
rect 3149 8132 3153 8188
rect 3089 8128 3153 8132
rect 6644 8188 6708 8192
rect 6644 8132 6648 8188
rect 6648 8132 6704 8188
rect 6704 8132 6708 8188
rect 6644 8128 6708 8132
rect 6724 8188 6788 8192
rect 6724 8132 6728 8188
rect 6728 8132 6784 8188
rect 6784 8132 6788 8188
rect 6724 8128 6788 8132
rect 6804 8188 6868 8192
rect 6804 8132 6808 8188
rect 6808 8132 6864 8188
rect 6864 8132 6868 8188
rect 6804 8128 6868 8132
rect 6884 8188 6948 8192
rect 6884 8132 6888 8188
rect 6888 8132 6944 8188
rect 6944 8132 6948 8188
rect 6884 8128 6948 8132
rect 10439 8188 10503 8192
rect 10439 8132 10443 8188
rect 10443 8132 10499 8188
rect 10499 8132 10503 8188
rect 10439 8128 10503 8132
rect 10519 8188 10583 8192
rect 10519 8132 10523 8188
rect 10523 8132 10579 8188
rect 10579 8132 10583 8188
rect 10519 8128 10583 8132
rect 10599 8188 10663 8192
rect 10599 8132 10603 8188
rect 10603 8132 10659 8188
rect 10659 8132 10663 8188
rect 10599 8128 10663 8132
rect 10679 8188 10743 8192
rect 10679 8132 10683 8188
rect 10683 8132 10739 8188
rect 10739 8132 10743 8188
rect 10679 8128 10743 8132
rect 14234 8188 14298 8192
rect 14234 8132 14238 8188
rect 14238 8132 14294 8188
rect 14294 8132 14298 8188
rect 14234 8128 14298 8132
rect 14314 8188 14378 8192
rect 14314 8132 14318 8188
rect 14318 8132 14374 8188
rect 14374 8132 14378 8188
rect 14314 8128 14378 8132
rect 14394 8188 14458 8192
rect 14394 8132 14398 8188
rect 14398 8132 14454 8188
rect 14454 8132 14458 8188
rect 14394 8128 14458 8132
rect 14474 8188 14538 8192
rect 14474 8132 14478 8188
rect 14478 8132 14534 8188
rect 14534 8132 14538 8188
rect 14474 8128 14538 8132
rect 3509 7644 3573 7648
rect 3509 7588 3513 7644
rect 3513 7588 3569 7644
rect 3569 7588 3573 7644
rect 3509 7584 3573 7588
rect 3589 7644 3653 7648
rect 3589 7588 3593 7644
rect 3593 7588 3649 7644
rect 3649 7588 3653 7644
rect 3589 7584 3653 7588
rect 3669 7644 3733 7648
rect 3669 7588 3673 7644
rect 3673 7588 3729 7644
rect 3729 7588 3733 7644
rect 3669 7584 3733 7588
rect 3749 7644 3813 7648
rect 3749 7588 3753 7644
rect 3753 7588 3809 7644
rect 3809 7588 3813 7644
rect 3749 7584 3813 7588
rect 7304 7644 7368 7648
rect 7304 7588 7308 7644
rect 7308 7588 7364 7644
rect 7364 7588 7368 7644
rect 7304 7584 7368 7588
rect 7384 7644 7448 7648
rect 7384 7588 7388 7644
rect 7388 7588 7444 7644
rect 7444 7588 7448 7644
rect 7384 7584 7448 7588
rect 7464 7644 7528 7648
rect 7464 7588 7468 7644
rect 7468 7588 7524 7644
rect 7524 7588 7528 7644
rect 7464 7584 7528 7588
rect 7544 7644 7608 7648
rect 7544 7588 7548 7644
rect 7548 7588 7604 7644
rect 7604 7588 7608 7644
rect 7544 7584 7608 7588
rect 11099 7644 11163 7648
rect 11099 7588 11103 7644
rect 11103 7588 11159 7644
rect 11159 7588 11163 7644
rect 11099 7584 11163 7588
rect 11179 7644 11243 7648
rect 11179 7588 11183 7644
rect 11183 7588 11239 7644
rect 11239 7588 11243 7644
rect 11179 7584 11243 7588
rect 11259 7644 11323 7648
rect 11259 7588 11263 7644
rect 11263 7588 11319 7644
rect 11319 7588 11323 7644
rect 11259 7584 11323 7588
rect 11339 7644 11403 7648
rect 11339 7588 11343 7644
rect 11343 7588 11399 7644
rect 11399 7588 11403 7644
rect 11339 7584 11403 7588
rect 14894 7644 14958 7648
rect 14894 7588 14898 7644
rect 14898 7588 14954 7644
rect 14954 7588 14958 7644
rect 14894 7584 14958 7588
rect 14974 7644 15038 7648
rect 14974 7588 14978 7644
rect 14978 7588 15034 7644
rect 15034 7588 15038 7644
rect 14974 7584 15038 7588
rect 15054 7644 15118 7648
rect 15054 7588 15058 7644
rect 15058 7588 15114 7644
rect 15114 7588 15118 7644
rect 15054 7584 15118 7588
rect 15134 7644 15198 7648
rect 15134 7588 15138 7644
rect 15138 7588 15194 7644
rect 15194 7588 15198 7644
rect 15134 7584 15198 7588
rect 2849 7100 2913 7104
rect 2849 7044 2853 7100
rect 2853 7044 2909 7100
rect 2909 7044 2913 7100
rect 2849 7040 2913 7044
rect 2929 7100 2993 7104
rect 2929 7044 2933 7100
rect 2933 7044 2989 7100
rect 2989 7044 2993 7100
rect 2929 7040 2993 7044
rect 3009 7100 3073 7104
rect 3009 7044 3013 7100
rect 3013 7044 3069 7100
rect 3069 7044 3073 7100
rect 3009 7040 3073 7044
rect 3089 7100 3153 7104
rect 3089 7044 3093 7100
rect 3093 7044 3149 7100
rect 3149 7044 3153 7100
rect 3089 7040 3153 7044
rect 6644 7100 6708 7104
rect 6644 7044 6648 7100
rect 6648 7044 6704 7100
rect 6704 7044 6708 7100
rect 6644 7040 6708 7044
rect 6724 7100 6788 7104
rect 6724 7044 6728 7100
rect 6728 7044 6784 7100
rect 6784 7044 6788 7100
rect 6724 7040 6788 7044
rect 6804 7100 6868 7104
rect 6804 7044 6808 7100
rect 6808 7044 6864 7100
rect 6864 7044 6868 7100
rect 6804 7040 6868 7044
rect 6884 7100 6948 7104
rect 6884 7044 6888 7100
rect 6888 7044 6944 7100
rect 6944 7044 6948 7100
rect 6884 7040 6948 7044
rect 10439 7100 10503 7104
rect 10439 7044 10443 7100
rect 10443 7044 10499 7100
rect 10499 7044 10503 7100
rect 10439 7040 10503 7044
rect 10519 7100 10583 7104
rect 10519 7044 10523 7100
rect 10523 7044 10579 7100
rect 10579 7044 10583 7100
rect 10519 7040 10583 7044
rect 10599 7100 10663 7104
rect 10599 7044 10603 7100
rect 10603 7044 10659 7100
rect 10659 7044 10663 7100
rect 10599 7040 10663 7044
rect 10679 7100 10743 7104
rect 10679 7044 10683 7100
rect 10683 7044 10739 7100
rect 10739 7044 10743 7100
rect 10679 7040 10743 7044
rect 14234 7100 14298 7104
rect 14234 7044 14238 7100
rect 14238 7044 14294 7100
rect 14294 7044 14298 7100
rect 14234 7040 14298 7044
rect 14314 7100 14378 7104
rect 14314 7044 14318 7100
rect 14318 7044 14374 7100
rect 14374 7044 14378 7100
rect 14314 7040 14378 7044
rect 14394 7100 14458 7104
rect 14394 7044 14398 7100
rect 14398 7044 14454 7100
rect 14454 7044 14458 7100
rect 14394 7040 14458 7044
rect 14474 7100 14538 7104
rect 14474 7044 14478 7100
rect 14478 7044 14534 7100
rect 14534 7044 14538 7100
rect 14474 7040 14538 7044
rect 3509 6556 3573 6560
rect 3509 6500 3513 6556
rect 3513 6500 3569 6556
rect 3569 6500 3573 6556
rect 3509 6496 3573 6500
rect 3589 6556 3653 6560
rect 3589 6500 3593 6556
rect 3593 6500 3649 6556
rect 3649 6500 3653 6556
rect 3589 6496 3653 6500
rect 3669 6556 3733 6560
rect 3669 6500 3673 6556
rect 3673 6500 3729 6556
rect 3729 6500 3733 6556
rect 3669 6496 3733 6500
rect 3749 6556 3813 6560
rect 3749 6500 3753 6556
rect 3753 6500 3809 6556
rect 3809 6500 3813 6556
rect 3749 6496 3813 6500
rect 7304 6556 7368 6560
rect 7304 6500 7308 6556
rect 7308 6500 7364 6556
rect 7364 6500 7368 6556
rect 7304 6496 7368 6500
rect 7384 6556 7448 6560
rect 7384 6500 7388 6556
rect 7388 6500 7444 6556
rect 7444 6500 7448 6556
rect 7384 6496 7448 6500
rect 7464 6556 7528 6560
rect 7464 6500 7468 6556
rect 7468 6500 7524 6556
rect 7524 6500 7528 6556
rect 7464 6496 7528 6500
rect 7544 6556 7608 6560
rect 7544 6500 7548 6556
rect 7548 6500 7604 6556
rect 7604 6500 7608 6556
rect 7544 6496 7608 6500
rect 11099 6556 11163 6560
rect 11099 6500 11103 6556
rect 11103 6500 11159 6556
rect 11159 6500 11163 6556
rect 11099 6496 11163 6500
rect 11179 6556 11243 6560
rect 11179 6500 11183 6556
rect 11183 6500 11239 6556
rect 11239 6500 11243 6556
rect 11179 6496 11243 6500
rect 11259 6556 11323 6560
rect 11259 6500 11263 6556
rect 11263 6500 11319 6556
rect 11319 6500 11323 6556
rect 11259 6496 11323 6500
rect 11339 6556 11403 6560
rect 11339 6500 11343 6556
rect 11343 6500 11399 6556
rect 11399 6500 11403 6556
rect 11339 6496 11403 6500
rect 14894 6556 14958 6560
rect 14894 6500 14898 6556
rect 14898 6500 14954 6556
rect 14954 6500 14958 6556
rect 14894 6496 14958 6500
rect 14974 6556 15038 6560
rect 14974 6500 14978 6556
rect 14978 6500 15034 6556
rect 15034 6500 15038 6556
rect 14974 6496 15038 6500
rect 15054 6556 15118 6560
rect 15054 6500 15058 6556
rect 15058 6500 15114 6556
rect 15114 6500 15118 6556
rect 15054 6496 15118 6500
rect 15134 6556 15198 6560
rect 15134 6500 15138 6556
rect 15138 6500 15194 6556
rect 15194 6500 15198 6556
rect 15134 6496 15198 6500
rect 2849 6012 2913 6016
rect 2849 5956 2853 6012
rect 2853 5956 2909 6012
rect 2909 5956 2913 6012
rect 2849 5952 2913 5956
rect 2929 6012 2993 6016
rect 2929 5956 2933 6012
rect 2933 5956 2989 6012
rect 2989 5956 2993 6012
rect 2929 5952 2993 5956
rect 3009 6012 3073 6016
rect 3009 5956 3013 6012
rect 3013 5956 3069 6012
rect 3069 5956 3073 6012
rect 3009 5952 3073 5956
rect 3089 6012 3153 6016
rect 3089 5956 3093 6012
rect 3093 5956 3149 6012
rect 3149 5956 3153 6012
rect 3089 5952 3153 5956
rect 6644 6012 6708 6016
rect 6644 5956 6648 6012
rect 6648 5956 6704 6012
rect 6704 5956 6708 6012
rect 6644 5952 6708 5956
rect 6724 6012 6788 6016
rect 6724 5956 6728 6012
rect 6728 5956 6784 6012
rect 6784 5956 6788 6012
rect 6724 5952 6788 5956
rect 6804 6012 6868 6016
rect 6804 5956 6808 6012
rect 6808 5956 6864 6012
rect 6864 5956 6868 6012
rect 6804 5952 6868 5956
rect 6884 6012 6948 6016
rect 6884 5956 6888 6012
rect 6888 5956 6944 6012
rect 6944 5956 6948 6012
rect 6884 5952 6948 5956
rect 10439 6012 10503 6016
rect 10439 5956 10443 6012
rect 10443 5956 10499 6012
rect 10499 5956 10503 6012
rect 10439 5952 10503 5956
rect 10519 6012 10583 6016
rect 10519 5956 10523 6012
rect 10523 5956 10579 6012
rect 10579 5956 10583 6012
rect 10519 5952 10583 5956
rect 10599 6012 10663 6016
rect 10599 5956 10603 6012
rect 10603 5956 10659 6012
rect 10659 5956 10663 6012
rect 10599 5952 10663 5956
rect 10679 6012 10743 6016
rect 10679 5956 10683 6012
rect 10683 5956 10739 6012
rect 10739 5956 10743 6012
rect 10679 5952 10743 5956
rect 14234 6012 14298 6016
rect 14234 5956 14238 6012
rect 14238 5956 14294 6012
rect 14294 5956 14298 6012
rect 14234 5952 14298 5956
rect 14314 6012 14378 6016
rect 14314 5956 14318 6012
rect 14318 5956 14374 6012
rect 14374 5956 14378 6012
rect 14314 5952 14378 5956
rect 14394 6012 14458 6016
rect 14394 5956 14398 6012
rect 14398 5956 14454 6012
rect 14454 5956 14458 6012
rect 14394 5952 14458 5956
rect 14474 6012 14538 6016
rect 14474 5956 14478 6012
rect 14478 5956 14534 6012
rect 14534 5956 14538 6012
rect 14474 5952 14538 5956
rect 3509 5468 3573 5472
rect 3509 5412 3513 5468
rect 3513 5412 3569 5468
rect 3569 5412 3573 5468
rect 3509 5408 3573 5412
rect 3589 5468 3653 5472
rect 3589 5412 3593 5468
rect 3593 5412 3649 5468
rect 3649 5412 3653 5468
rect 3589 5408 3653 5412
rect 3669 5468 3733 5472
rect 3669 5412 3673 5468
rect 3673 5412 3729 5468
rect 3729 5412 3733 5468
rect 3669 5408 3733 5412
rect 3749 5468 3813 5472
rect 3749 5412 3753 5468
rect 3753 5412 3809 5468
rect 3809 5412 3813 5468
rect 3749 5408 3813 5412
rect 7304 5468 7368 5472
rect 7304 5412 7308 5468
rect 7308 5412 7364 5468
rect 7364 5412 7368 5468
rect 7304 5408 7368 5412
rect 7384 5468 7448 5472
rect 7384 5412 7388 5468
rect 7388 5412 7444 5468
rect 7444 5412 7448 5468
rect 7384 5408 7448 5412
rect 7464 5468 7528 5472
rect 7464 5412 7468 5468
rect 7468 5412 7524 5468
rect 7524 5412 7528 5468
rect 7464 5408 7528 5412
rect 7544 5468 7608 5472
rect 7544 5412 7548 5468
rect 7548 5412 7604 5468
rect 7604 5412 7608 5468
rect 7544 5408 7608 5412
rect 11099 5468 11163 5472
rect 11099 5412 11103 5468
rect 11103 5412 11159 5468
rect 11159 5412 11163 5468
rect 11099 5408 11163 5412
rect 11179 5468 11243 5472
rect 11179 5412 11183 5468
rect 11183 5412 11239 5468
rect 11239 5412 11243 5468
rect 11179 5408 11243 5412
rect 11259 5468 11323 5472
rect 11259 5412 11263 5468
rect 11263 5412 11319 5468
rect 11319 5412 11323 5468
rect 11259 5408 11323 5412
rect 11339 5468 11403 5472
rect 11339 5412 11343 5468
rect 11343 5412 11399 5468
rect 11399 5412 11403 5468
rect 11339 5408 11403 5412
rect 14894 5468 14958 5472
rect 14894 5412 14898 5468
rect 14898 5412 14954 5468
rect 14954 5412 14958 5468
rect 14894 5408 14958 5412
rect 14974 5468 15038 5472
rect 14974 5412 14978 5468
rect 14978 5412 15034 5468
rect 15034 5412 15038 5468
rect 14974 5408 15038 5412
rect 15054 5468 15118 5472
rect 15054 5412 15058 5468
rect 15058 5412 15114 5468
rect 15114 5412 15118 5468
rect 15054 5408 15118 5412
rect 15134 5468 15198 5472
rect 15134 5412 15138 5468
rect 15138 5412 15194 5468
rect 15194 5412 15198 5468
rect 15134 5408 15198 5412
rect 2849 4924 2913 4928
rect 2849 4868 2853 4924
rect 2853 4868 2909 4924
rect 2909 4868 2913 4924
rect 2849 4864 2913 4868
rect 2929 4924 2993 4928
rect 2929 4868 2933 4924
rect 2933 4868 2989 4924
rect 2989 4868 2993 4924
rect 2929 4864 2993 4868
rect 3009 4924 3073 4928
rect 3009 4868 3013 4924
rect 3013 4868 3069 4924
rect 3069 4868 3073 4924
rect 3009 4864 3073 4868
rect 3089 4924 3153 4928
rect 3089 4868 3093 4924
rect 3093 4868 3149 4924
rect 3149 4868 3153 4924
rect 3089 4864 3153 4868
rect 6644 4924 6708 4928
rect 6644 4868 6648 4924
rect 6648 4868 6704 4924
rect 6704 4868 6708 4924
rect 6644 4864 6708 4868
rect 6724 4924 6788 4928
rect 6724 4868 6728 4924
rect 6728 4868 6784 4924
rect 6784 4868 6788 4924
rect 6724 4864 6788 4868
rect 6804 4924 6868 4928
rect 6804 4868 6808 4924
rect 6808 4868 6864 4924
rect 6864 4868 6868 4924
rect 6804 4864 6868 4868
rect 6884 4924 6948 4928
rect 6884 4868 6888 4924
rect 6888 4868 6944 4924
rect 6944 4868 6948 4924
rect 6884 4864 6948 4868
rect 10439 4924 10503 4928
rect 10439 4868 10443 4924
rect 10443 4868 10499 4924
rect 10499 4868 10503 4924
rect 10439 4864 10503 4868
rect 10519 4924 10583 4928
rect 10519 4868 10523 4924
rect 10523 4868 10579 4924
rect 10579 4868 10583 4924
rect 10519 4864 10583 4868
rect 10599 4924 10663 4928
rect 10599 4868 10603 4924
rect 10603 4868 10659 4924
rect 10659 4868 10663 4924
rect 10599 4864 10663 4868
rect 10679 4924 10743 4928
rect 10679 4868 10683 4924
rect 10683 4868 10739 4924
rect 10739 4868 10743 4924
rect 10679 4864 10743 4868
rect 14234 4924 14298 4928
rect 14234 4868 14238 4924
rect 14238 4868 14294 4924
rect 14294 4868 14298 4924
rect 14234 4864 14298 4868
rect 14314 4924 14378 4928
rect 14314 4868 14318 4924
rect 14318 4868 14374 4924
rect 14374 4868 14378 4924
rect 14314 4864 14378 4868
rect 14394 4924 14458 4928
rect 14394 4868 14398 4924
rect 14398 4868 14454 4924
rect 14454 4868 14458 4924
rect 14394 4864 14458 4868
rect 14474 4924 14538 4928
rect 14474 4868 14478 4924
rect 14478 4868 14534 4924
rect 14534 4868 14538 4924
rect 14474 4864 14538 4868
rect 3509 4380 3573 4384
rect 3509 4324 3513 4380
rect 3513 4324 3569 4380
rect 3569 4324 3573 4380
rect 3509 4320 3573 4324
rect 3589 4380 3653 4384
rect 3589 4324 3593 4380
rect 3593 4324 3649 4380
rect 3649 4324 3653 4380
rect 3589 4320 3653 4324
rect 3669 4380 3733 4384
rect 3669 4324 3673 4380
rect 3673 4324 3729 4380
rect 3729 4324 3733 4380
rect 3669 4320 3733 4324
rect 3749 4380 3813 4384
rect 3749 4324 3753 4380
rect 3753 4324 3809 4380
rect 3809 4324 3813 4380
rect 3749 4320 3813 4324
rect 7304 4380 7368 4384
rect 7304 4324 7308 4380
rect 7308 4324 7364 4380
rect 7364 4324 7368 4380
rect 7304 4320 7368 4324
rect 7384 4380 7448 4384
rect 7384 4324 7388 4380
rect 7388 4324 7444 4380
rect 7444 4324 7448 4380
rect 7384 4320 7448 4324
rect 7464 4380 7528 4384
rect 7464 4324 7468 4380
rect 7468 4324 7524 4380
rect 7524 4324 7528 4380
rect 7464 4320 7528 4324
rect 7544 4380 7608 4384
rect 7544 4324 7548 4380
rect 7548 4324 7604 4380
rect 7604 4324 7608 4380
rect 7544 4320 7608 4324
rect 11099 4380 11163 4384
rect 11099 4324 11103 4380
rect 11103 4324 11159 4380
rect 11159 4324 11163 4380
rect 11099 4320 11163 4324
rect 11179 4380 11243 4384
rect 11179 4324 11183 4380
rect 11183 4324 11239 4380
rect 11239 4324 11243 4380
rect 11179 4320 11243 4324
rect 11259 4380 11323 4384
rect 11259 4324 11263 4380
rect 11263 4324 11319 4380
rect 11319 4324 11323 4380
rect 11259 4320 11323 4324
rect 11339 4380 11403 4384
rect 11339 4324 11343 4380
rect 11343 4324 11399 4380
rect 11399 4324 11403 4380
rect 11339 4320 11403 4324
rect 14894 4380 14958 4384
rect 14894 4324 14898 4380
rect 14898 4324 14954 4380
rect 14954 4324 14958 4380
rect 14894 4320 14958 4324
rect 14974 4380 15038 4384
rect 14974 4324 14978 4380
rect 14978 4324 15034 4380
rect 15034 4324 15038 4380
rect 14974 4320 15038 4324
rect 15054 4380 15118 4384
rect 15054 4324 15058 4380
rect 15058 4324 15114 4380
rect 15114 4324 15118 4380
rect 15054 4320 15118 4324
rect 15134 4380 15198 4384
rect 15134 4324 15138 4380
rect 15138 4324 15194 4380
rect 15194 4324 15198 4380
rect 15134 4320 15198 4324
rect 2849 3836 2913 3840
rect 2849 3780 2853 3836
rect 2853 3780 2909 3836
rect 2909 3780 2913 3836
rect 2849 3776 2913 3780
rect 2929 3836 2993 3840
rect 2929 3780 2933 3836
rect 2933 3780 2989 3836
rect 2989 3780 2993 3836
rect 2929 3776 2993 3780
rect 3009 3836 3073 3840
rect 3009 3780 3013 3836
rect 3013 3780 3069 3836
rect 3069 3780 3073 3836
rect 3009 3776 3073 3780
rect 3089 3836 3153 3840
rect 3089 3780 3093 3836
rect 3093 3780 3149 3836
rect 3149 3780 3153 3836
rect 3089 3776 3153 3780
rect 6644 3836 6708 3840
rect 6644 3780 6648 3836
rect 6648 3780 6704 3836
rect 6704 3780 6708 3836
rect 6644 3776 6708 3780
rect 6724 3836 6788 3840
rect 6724 3780 6728 3836
rect 6728 3780 6784 3836
rect 6784 3780 6788 3836
rect 6724 3776 6788 3780
rect 6804 3836 6868 3840
rect 6804 3780 6808 3836
rect 6808 3780 6864 3836
rect 6864 3780 6868 3836
rect 6804 3776 6868 3780
rect 6884 3836 6948 3840
rect 6884 3780 6888 3836
rect 6888 3780 6944 3836
rect 6944 3780 6948 3836
rect 6884 3776 6948 3780
rect 10439 3836 10503 3840
rect 10439 3780 10443 3836
rect 10443 3780 10499 3836
rect 10499 3780 10503 3836
rect 10439 3776 10503 3780
rect 10519 3836 10583 3840
rect 10519 3780 10523 3836
rect 10523 3780 10579 3836
rect 10579 3780 10583 3836
rect 10519 3776 10583 3780
rect 10599 3836 10663 3840
rect 10599 3780 10603 3836
rect 10603 3780 10659 3836
rect 10659 3780 10663 3836
rect 10599 3776 10663 3780
rect 10679 3836 10743 3840
rect 10679 3780 10683 3836
rect 10683 3780 10739 3836
rect 10739 3780 10743 3836
rect 10679 3776 10743 3780
rect 14234 3836 14298 3840
rect 14234 3780 14238 3836
rect 14238 3780 14294 3836
rect 14294 3780 14298 3836
rect 14234 3776 14298 3780
rect 14314 3836 14378 3840
rect 14314 3780 14318 3836
rect 14318 3780 14374 3836
rect 14374 3780 14378 3836
rect 14314 3776 14378 3780
rect 14394 3836 14458 3840
rect 14394 3780 14398 3836
rect 14398 3780 14454 3836
rect 14454 3780 14458 3836
rect 14394 3776 14458 3780
rect 14474 3836 14538 3840
rect 14474 3780 14478 3836
rect 14478 3780 14534 3836
rect 14534 3780 14538 3836
rect 14474 3776 14538 3780
rect 3509 3292 3573 3296
rect 3509 3236 3513 3292
rect 3513 3236 3569 3292
rect 3569 3236 3573 3292
rect 3509 3232 3573 3236
rect 3589 3292 3653 3296
rect 3589 3236 3593 3292
rect 3593 3236 3649 3292
rect 3649 3236 3653 3292
rect 3589 3232 3653 3236
rect 3669 3292 3733 3296
rect 3669 3236 3673 3292
rect 3673 3236 3729 3292
rect 3729 3236 3733 3292
rect 3669 3232 3733 3236
rect 3749 3292 3813 3296
rect 3749 3236 3753 3292
rect 3753 3236 3809 3292
rect 3809 3236 3813 3292
rect 3749 3232 3813 3236
rect 7304 3292 7368 3296
rect 7304 3236 7308 3292
rect 7308 3236 7364 3292
rect 7364 3236 7368 3292
rect 7304 3232 7368 3236
rect 7384 3292 7448 3296
rect 7384 3236 7388 3292
rect 7388 3236 7444 3292
rect 7444 3236 7448 3292
rect 7384 3232 7448 3236
rect 7464 3292 7528 3296
rect 7464 3236 7468 3292
rect 7468 3236 7524 3292
rect 7524 3236 7528 3292
rect 7464 3232 7528 3236
rect 7544 3292 7608 3296
rect 7544 3236 7548 3292
rect 7548 3236 7604 3292
rect 7604 3236 7608 3292
rect 7544 3232 7608 3236
rect 11099 3292 11163 3296
rect 11099 3236 11103 3292
rect 11103 3236 11159 3292
rect 11159 3236 11163 3292
rect 11099 3232 11163 3236
rect 11179 3292 11243 3296
rect 11179 3236 11183 3292
rect 11183 3236 11239 3292
rect 11239 3236 11243 3292
rect 11179 3232 11243 3236
rect 11259 3292 11323 3296
rect 11259 3236 11263 3292
rect 11263 3236 11319 3292
rect 11319 3236 11323 3292
rect 11259 3232 11323 3236
rect 11339 3292 11403 3296
rect 11339 3236 11343 3292
rect 11343 3236 11399 3292
rect 11399 3236 11403 3292
rect 11339 3232 11403 3236
rect 14894 3292 14958 3296
rect 14894 3236 14898 3292
rect 14898 3236 14954 3292
rect 14954 3236 14958 3292
rect 14894 3232 14958 3236
rect 14974 3292 15038 3296
rect 14974 3236 14978 3292
rect 14978 3236 15034 3292
rect 15034 3236 15038 3292
rect 14974 3232 15038 3236
rect 15054 3292 15118 3296
rect 15054 3236 15058 3292
rect 15058 3236 15114 3292
rect 15114 3236 15118 3292
rect 15054 3232 15118 3236
rect 15134 3292 15198 3296
rect 15134 3236 15138 3292
rect 15138 3236 15194 3292
rect 15194 3236 15198 3292
rect 15134 3232 15198 3236
rect 2849 2748 2913 2752
rect 2849 2692 2853 2748
rect 2853 2692 2909 2748
rect 2909 2692 2913 2748
rect 2849 2688 2913 2692
rect 2929 2748 2993 2752
rect 2929 2692 2933 2748
rect 2933 2692 2989 2748
rect 2989 2692 2993 2748
rect 2929 2688 2993 2692
rect 3009 2748 3073 2752
rect 3009 2692 3013 2748
rect 3013 2692 3069 2748
rect 3069 2692 3073 2748
rect 3009 2688 3073 2692
rect 3089 2748 3153 2752
rect 3089 2692 3093 2748
rect 3093 2692 3149 2748
rect 3149 2692 3153 2748
rect 3089 2688 3153 2692
rect 6644 2748 6708 2752
rect 6644 2692 6648 2748
rect 6648 2692 6704 2748
rect 6704 2692 6708 2748
rect 6644 2688 6708 2692
rect 6724 2748 6788 2752
rect 6724 2692 6728 2748
rect 6728 2692 6784 2748
rect 6784 2692 6788 2748
rect 6724 2688 6788 2692
rect 6804 2748 6868 2752
rect 6804 2692 6808 2748
rect 6808 2692 6864 2748
rect 6864 2692 6868 2748
rect 6804 2688 6868 2692
rect 6884 2748 6948 2752
rect 6884 2692 6888 2748
rect 6888 2692 6944 2748
rect 6944 2692 6948 2748
rect 6884 2688 6948 2692
rect 10439 2748 10503 2752
rect 10439 2692 10443 2748
rect 10443 2692 10499 2748
rect 10499 2692 10503 2748
rect 10439 2688 10503 2692
rect 10519 2748 10583 2752
rect 10519 2692 10523 2748
rect 10523 2692 10579 2748
rect 10579 2692 10583 2748
rect 10519 2688 10583 2692
rect 10599 2748 10663 2752
rect 10599 2692 10603 2748
rect 10603 2692 10659 2748
rect 10659 2692 10663 2748
rect 10599 2688 10663 2692
rect 10679 2748 10743 2752
rect 10679 2692 10683 2748
rect 10683 2692 10739 2748
rect 10739 2692 10743 2748
rect 10679 2688 10743 2692
rect 14234 2748 14298 2752
rect 14234 2692 14238 2748
rect 14238 2692 14294 2748
rect 14294 2692 14298 2748
rect 14234 2688 14298 2692
rect 14314 2748 14378 2752
rect 14314 2692 14318 2748
rect 14318 2692 14374 2748
rect 14374 2692 14378 2748
rect 14314 2688 14378 2692
rect 14394 2748 14458 2752
rect 14394 2692 14398 2748
rect 14398 2692 14454 2748
rect 14454 2692 14458 2748
rect 14394 2688 14458 2692
rect 14474 2748 14538 2752
rect 14474 2692 14478 2748
rect 14478 2692 14534 2748
rect 14534 2692 14538 2748
rect 14474 2688 14538 2692
rect 3509 2204 3573 2208
rect 3509 2148 3513 2204
rect 3513 2148 3569 2204
rect 3569 2148 3573 2204
rect 3509 2144 3573 2148
rect 3589 2204 3653 2208
rect 3589 2148 3593 2204
rect 3593 2148 3649 2204
rect 3649 2148 3653 2204
rect 3589 2144 3653 2148
rect 3669 2204 3733 2208
rect 3669 2148 3673 2204
rect 3673 2148 3729 2204
rect 3729 2148 3733 2204
rect 3669 2144 3733 2148
rect 3749 2204 3813 2208
rect 3749 2148 3753 2204
rect 3753 2148 3809 2204
rect 3809 2148 3813 2204
rect 3749 2144 3813 2148
rect 7304 2204 7368 2208
rect 7304 2148 7308 2204
rect 7308 2148 7364 2204
rect 7364 2148 7368 2204
rect 7304 2144 7368 2148
rect 7384 2204 7448 2208
rect 7384 2148 7388 2204
rect 7388 2148 7444 2204
rect 7444 2148 7448 2204
rect 7384 2144 7448 2148
rect 7464 2204 7528 2208
rect 7464 2148 7468 2204
rect 7468 2148 7524 2204
rect 7524 2148 7528 2204
rect 7464 2144 7528 2148
rect 7544 2204 7608 2208
rect 7544 2148 7548 2204
rect 7548 2148 7604 2204
rect 7604 2148 7608 2204
rect 7544 2144 7608 2148
rect 11099 2204 11163 2208
rect 11099 2148 11103 2204
rect 11103 2148 11159 2204
rect 11159 2148 11163 2204
rect 11099 2144 11163 2148
rect 11179 2204 11243 2208
rect 11179 2148 11183 2204
rect 11183 2148 11239 2204
rect 11239 2148 11243 2204
rect 11179 2144 11243 2148
rect 11259 2204 11323 2208
rect 11259 2148 11263 2204
rect 11263 2148 11319 2204
rect 11319 2148 11323 2204
rect 11259 2144 11323 2148
rect 11339 2204 11403 2208
rect 11339 2148 11343 2204
rect 11343 2148 11399 2204
rect 11399 2148 11403 2204
rect 11339 2144 11403 2148
rect 14894 2204 14958 2208
rect 14894 2148 14898 2204
rect 14898 2148 14954 2204
rect 14954 2148 14958 2204
rect 14894 2144 14958 2148
rect 14974 2204 15038 2208
rect 14974 2148 14978 2204
rect 14978 2148 15034 2204
rect 15034 2148 15038 2204
rect 14974 2144 15038 2148
rect 15054 2204 15118 2208
rect 15054 2148 15058 2204
rect 15058 2148 15114 2204
rect 15114 2148 15118 2204
rect 15054 2144 15118 2148
rect 15134 2204 15198 2208
rect 15134 2148 15138 2204
rect 15138 2148 15194 2204
rect 15194 2148 15198 2204
rect 15134 2144 15198 2148
<< metal4 >>
rect 2841 16896 3161 16912
rect 2841 16832 2849 16896
rect 2913 16832 2929 16896
rect 2993 16832 3009 16896
rect 3073 16832 3089 16896
rect 3153 16832 3161 16896
rect 2841 15808 3161 16832
rect 2841 15744 2849 15808
rect 2913 15744 2929 15808
rect 2993 15744 3009 15808
rect 3073 15744 3089 15808
rect 3153 15744 3161 15808
rect 2841 15146 3161 15744
rect 2841 14910 2883 15146
rect 3119 14910 3161 15146
rect 2841 14720 3161 14910
rect 2841 14656 2849 14720
rect 2913 14656 2929 14720
rect 2993 14656 3009 14720
rect 3073 14656 3089 14720
rect 3153 14656 3161 14720
rect 2841 13632 3161 14656
rect 2841 13568 2849 13632
rect 2913 13568 2929 13632
rect 2993 13568 3009 13632
rect 3073 13568 3089 13632
rect 3153 13568 3161 13632
rect 2841 12544 3161 13568
rect 2841 12480 2849 12544
rect 2913 12480 2929 12544
rect 2993 12480 3009 12544
rect 3073 12480 3089 12544
rect 3153 12480 3161 12544
rect 2841 11474 3161 12480
rect 2841 11456 2883 11474
rect 3119 11456 3161 11474
rect 2841 11392 2849 11456
rect 3153 11392 3161 11456
rect 2841 11238 2883 11392
rect 3119 11238 3161 11392
rect 2841 10368 3161 11238
rect 2841 10304 2849 10368
rect 2913 10304 2929 10368
rect 2993 10304 3009 10368
rect 3073 10304 3089 10368
rect 3153 10304 3161 10368
rect 2841 9280 3161 10304
rect 2841 9216 2849 9280
rect 2913 9216 2929 9280
rect 2993 9216 3009 9280
rect 3073 9216 3089 9280
rect 3153 9216 3161 9280
rect 2841 8192 3161 9216
rect 2841 8128 2849 8192
rect 2913 8128 2929 8192
rect 2993 8128 3009 8192
rect 3073 8128 3089 8192
rect 3153 8128 3161 8192
rect 2841 7802 3161 8128
rect 2841 7566 2883 7802
rect 3119 7566 3161 7802
rect 2841 7104 3161 7566
rect 2841 7040 2849 7104
rect 2913 7040 2929 7104
rect 2993 7040 3009 7104
rect 3073 7040 3089 7104
rect 3153 7040 3161 7104
rect 2841 6016 3161 7040
rect 2841 5952 2849 6016
rect 2913 5952 2929 6016
rect 2993 5952 3009 6016
rect 3073 5952 3089 6016
rect 3153 5952 3161 6016
rect 2841 4928 3161 5952
rect 2841 4864 2849 4928
rect 2913 4864 2929 4928
rect 2993 4864 3009 4928
rect 3073 4864 3089 4928
rect 3153 4864 3161 4928
rect 2841 4130 3161 4864
rect 2841 3894 2883 4130
rect 3119 3894 3161 4130
rect 2841 3840 3161 3894
rect 2841 3776 2849 3840
rect 2913 3776 2929 3840
rect 2993 3776 3009 3840
rect 3073 3776 3089 3840
rect 3153 3776 3161 3840
rect 2841 2752 3161 3776
rect 2841 2688 2849 2752
rect 2913 2688 2929 2752
rect 2993 2688 3009 2752
rect 3073 2688 3089 2752
rect 3153 2688 3161 2752
rect 2841 2128 3161 2688
rect 3501 16352 3821 16912
rect 3501 16288 3509 16352
rect 3573 16288 3589 16352
rect 3653 16288 3669 16352
rect 3733 16288 3749 16352
rect 3813 16288 3821 16352
rect 3501 15806 3821 16288
rect 3501 15570 3543 15806
rect 3779 15570 3821 15806
rect 3501 15264 3821 15570
rect 3501 15200 3509 15264
rect 3573 15200 3589 15264
rect 3653 15200 3669 15264
rect 3733 15200 3749 15264
rect 3813 15200 3821 15264
rect 3501 14176 3821 15200
rect 3501 14112 3509 14176
rect 3573 14112 3589 14176
rect 3653 14112 3669 14176
rect 3733 14112 3749 14176
rect 3813 14112 3821 14176
rect 3501 13088 3821 14112
rect 3501 13024 3509 13088
rect 3573 13024 3589 13088
rect 3653 13024 3669 13088
rect 3733 13024 3749 13088
rect 3813 13024 3821 13088
rect 3501 12134 3821 13024
rect 3501 12000 3543 12134
rect 3779 12000 3821 12134
rect 3501 11936 3509 12000
rect 3813 11936 3821 12000
rect 3501 11898 3543 11936
rect 3779 11898 3821 11936
rect 3501 10912 3821 11898
rect 3501 10848 3509 10912
rect 3573 10848 3589 10912
rect 3653 10848 3669 10912
rect 3733 10848 3749 10912
rect 3813 10848 3821 10912
rect 3501 9824 3821 10848
rect 3501 9760 3509 9824
rect 3573 9760 3589 9824
rect 3653 9760 3669 9824
rect 3733 9760 3749 9824
rect 3813 9760 3821 9824
rect 3501 8736 3821 9760
rect 3501 8672 3509 8736
rect 3573 8672 3589 8736
rect 3653 8672 3669 8736
rect 3733 8672 3749 8736
rect 3813 8672 3821 8736
rect 3501 8462 3821 8672
rect 3501 8226 3543 8462
rect 3779 8226 3821 8462
rect 3501 7648 3821 8226
rect 3501 7584 3509 7648
rect 3573 7584 3589 7648
rect 3653 7584 3669 7648
rect 3733 7584 3749 7648
rect 3813 7584 3821 7648
rect 3501 6560 3821 7584
rect 3501 6496 3509 6560
rect 3573 6496 3589 6560
rect 3653 6496 3669 6560
rect 3733 6496 3749 6560
rect 3813 6496 3821 6560
rect 3501 5472 3821 6496
rect 3501 5408 3509 5472
rect 3573 5408 3589 5472
rect 3653 5408 3669 5472
rect 3733 5408 3749 5472
rect 3813 5408 3821 5472
rect 3501 4790 3821 5408
rect 3501 4554 3543 4790
rect 3779 4554 3821 4790
rect 3501 4384 3821 4554
rect 3501 4320 3509 4384
rect 3573 4320 3589 4384
rect 3653 4320 3669 4384
rect 3733 4320 3749 4384
rect 3813 4320 3821 4384
rect 3501 3296 3821 4320
rect 3501 3232 3509 3296
rect 3573 3232 3589 3296
rect 3653 3232 3669 3296
rect 3733 3232 3749 3296
rect 3813 3232 3821 3296
rect 3501 2208 3821 3232
rect 3501 2144 3509 2208
rect 3573 2144 3589 2208
rect 3653 2144 3669 2208
rect 3733 2144 3749 2208
rect 3813 2144 3821 2208
rect 3501 2128 3821 2144
rect 6636 16896 6956 16912
rect 6636 16832 6644 16896
rect 6708 16832 6724 16896
rect 6788 16832 6804 16896
rect 6868 16832 6884 16896
rect 6948 16832 6956 16896
rect 6636 15808 6956 16832
rect 6636 15744 6644 15808
rect 6708 15744 6724 15808
rect 6788 15744 6804 15808
rect 6868 15744 6884 15808
rect 6948 15744 6956 15808
rect 6636 15146 6956 15744
rect 6636 14910 6678 15146
rect 6914 14910 6956 15146
rect 6636 14720 6956 14910
rect 6636 14656 6644 14720
rect 6708 14656 6724 14720
rect 6788 14656 6804 14720
rect 6868 14656 6884 14720
rect 6948 14656 6956 14720
rect 6636 13632 6956 14656
rect 6636 13568 6644 13632
rect 6708 13568 6724 13632
rect 6788 13568 6804 13632
rect 6868 13568 6884 13632
rect 6948 13568 6956 13632
rect 6636 12544 6956 13568
rect 6636 12480 6644 12544
rect 6708 12480 6724 12544
rect 6788 12480 6804 12544
rect 6868 12480 6884 12544
rect 6948 12480 6956 12544
rect 6636 11474 6956 12480
rect 6636 11456 6678 11474
rect 6914 11456 6956 11474
rect 6636 11392 6644 11456
rect 6948 11392 6956 11456
rect 6636 11238 6678 11392
rect 6914 11238 6956 11392
rect 6636 10368 6956 11238
rect 6636 10304 6644 10368
rect 6708 10304 6724 10368
rect 6788 10304 6804 10368
rect 6868 10304 6884 10368
rect 6948 10304 6956 10368
rect 6636 9280 6956 10304
rect 6636 9216 6644 9280
rect 6708 9216 6724 9280
rect 6788 9216 6804 9280
rect 6868 9216 6884 9280
rect 6948 9216 6956 9280
rect 6636 8192 6956 9216
rect 6636 8128 6644 8192
rect 6708 8128 6724 8192
rect 6788 8128 6804 8192
rect 6868 8128 6884 8192
rect 6948 8128 6956 8192
rect 6636 7802 6956 8128
rect 6636 7566 6678 7802
rect 6914 7566 6956 7802
rect 6636 7104 6956 7566
rect 6636 7040 6644 7104
rect 6708 7040 6724 7104
rect 6788 7040 6804 7104
rect 6868 7040 6884 7104
rect 6948 7040 6956 7104
rect 6636 6016 6956 7040
rect 6636 5952 6644 6016
rect 6708 5952 6724 6016
rect 6788 5952 6804 6016
rect 6868 5952 6884 6016
rect 6948 5952 6956 6016
rect 6636 4928 6956 5952
rect 6636 4864 6644 4928
rect 6708 4864 6724 4928
rect 6788 4864 6804 4928
rect 6868 4864 6884 4928
rect 6948 4864 6956 4928
rect 6636 4130 6956 4864
rect 6636 3894 6678 4130
rect 6914 3894 6956 4130
rect 6636 3840 6956 3894
rect 6636 3776 6644 3840
rect 6708 3776 6724 3840
rect 6788 3776 6804 3840
rect 6868 3776 6884 3840
rect 6948 3776 6956 3840
rect 6636 2752 6956 3776
rect 6636 2688 6644 2752
rect 6708 2688 6724 2752
rect 6788 2688 6804 2752
rect 6868 2688 6884 2752
rect 6948 2688 6956 2752
rect 6636 2128 6956 2688
rect 7296 16352 7616 16912
rect 7296 16288 7304 16352
rect 7368 16288 7384 16352
rect 7448 16288 7464 16352
rect 7528 16288 7544 16352
rect 7608 16288 7616 16352
rect 7296 15806 7616 16288
rect 7296 15570 7338 15806
rect 7574 15570 7616 15806
rect 7296 15264 7616 15570
rect 7296 15200 7304 15264
rect 7368 15200 7384 15264
rect 7448 15200 7464 15264
rect 7528 15200 7544 15264
rect 7608 15200 7616 15264
rect 7296 14176 7616 15200
rect 7296 14112 7304 14176
rect 7368 14112 7384 14176
rect 7448 14112 7464 14176
rect 7528 14112 7544 14176
rect 7608 14112 7616 14176
rect 7296 13088 7616 14112
rect 7296 13024 7304 13088
rect 7368 13024 7384 13088
rect 7448 13024 7464 13088
rect 7528 13024 7544 13088
rect 7608 13024 7616 13088
rect 7296 12134 7616 13024
rect 7296 12000 7338 12134
rect 7574 12000 7616 12134
rect 7296 11936 7304 12000
rect 7608 11936 7616 12000
rect 7296 11898 7338 11936
rect 7574 11898 7616 11936
rect 7296 10912 7616 11898
rect 7296 10848 7304 10912
rect 7368 10848 7384 10912
rect 7448 10848 7464 10912
rect 7528 10848 7544 10912
rect 7608 10848 7616 10912
rect 7296 9824 7616 10848
rect 7296 9760 7304 9824
rect 7368 9760 7384 9824
rect 7448 9760 7464 9824
rect 7528 9760 7544 9824
rect 7608 9760 7616 9824
rect 7296 8736 7616 9760
rect 7296 8672 7304 8736
rect 7368 8672 7384 8736
rect 7448 8672 7464 8736
rect 7528 8672 7544 8736
rect 7608 8672 7616 8736
rect 7296 8462 7616 8672
rect 7296 8226 7338 8462
rect 7574 8226 7616 8462
rect 7296 7648 7616 8226
rect 7296 7584 7304 7648
rect 7368 7584 7384 7648
rect 7448 7584 7464 7648
rect 7528 7584 7544 7648
rect 7608 7584 7616 7648
rect 7296 6560 7616 7584
rect 7296 6496 7304 6560
rect 7368 6496 7384 6560
rect 7448 6496 7464 6560
rect 7528 6496 7544 6560
rect 7608 6496 7616 6560
rect 7296 5472 7616 6496
rect 7296 5408 7304 5472
rect 7368 5408 7384 5472
rect 7448 5408 7464 5472
rect 7528 5408 7544 5472
rect 7608 5408 7616 5472
rect 7296 4790 7616 5408
rect 7296 4554 7338 4790
rect 7574 4554 7616 4790
rect 7296 4384 7616 4554
rect 7296 4320 7304 4384
rect 7368 4320 7384 4384
rect 7448 4320 7464 4384
rect 7528 4320 7544 4384
rect 7608 4320 7616 4384
rect 7296 3296 7616 4320
rect 7296 3232 7304 3296
rect 7368 3232 7384 3296
rect 7448 3232 7464 3296
rect 7528 3232 7544 3296
rect 7608 3232 7616 3296
rect 7296 2208 7616 3232
rect 7296 2144 7304 2208
rect 7368 2144 7384 2208
rect 7448 2144 7464 2208
rect 7528 2144 7544 2208
rect 7608 2144 7616 2208
rect 7296 2128 7616 2144
rect 10431 16896 10751 16912
rect 10431 16832 10439 16896
rect 10503 16832 10519 16896
rect 10583 16832 10599 16896
rect 10663 16832 10679 16896
rect 10743 16832 10751 16896
rect 10431 15808 10751 16832
rect 10431 15744 10439 15808
rect 10503 15744 10519 15808
rect 10583 15744 10599 15808
rect 10663 15744 10679 15808
rect 10743 15744 10751 15808
rect 10431 15146 10751 15744
rect 10431 14910 10473 15146
rect 10709 14910 10751 15146
rect 10431 14720 10751 14910
rect 10431 14656 10439 14720
rect 10503 14656 10519 14720
rect 10583 14656 10599 14720
rect 10663 14656 10679 14720
rect 10743 14656 10751 14720
rect 10431 13632 10751 14656
rect 10431 13568 10439 13632
rect 10503 13568 10519 13632
rect 10583 13568 10599 13632
rect 10663 13568 10679 13632
rect 10743 13568 10751 13632
rect 10431 12544 10751 13568
rect 10431 12480 10439 12544
rect 10503 12480 10519 12544
rect 10583 12480 10599 12544
rect 10663 12480 10679 12544
rect 10743 12480 10751 12544
rect 10431 11474 10751 12480
rect 10431 11456 10473 11474
rect 10709 11456 10751 11474
rect 10431 11392 10439 11456
rect 10743 11392 10751 11456
rect 10431 11238 10473 11392
rect 10709 11238 10751 11392
rect 10431 10368 10751 11238
rect 10431 10304 10439 10368
rect 10503 10304 10519 10368
rect 10583 10304 10599 10368
rect 10663 10304 10679 10368
rect 10743 10304 10751 10368
rect 10431 9280 10751 10304
rect 10431 9216 10439 9280
rect 10503 9216 10519 9280
rect 10583 9216 10599 9280
rect 10663 9216 10679 9280
rect 10743 9216 10751 9280
rect 10431 8192 10751 9216
rect 10431 8128 10439 8192
rect 10503 8128 10519 8192
rect 10583 8128 10599 8192
rect 10663 8128 10679 8192
rect 10743 8128 10751 8192
rect 10431 7802 10751 8128
rect 10431 7566 10473 7802
rect 10709 7566 10751 7802
rect 10431 7104 10751 7566
rect 10431 7040 10439 7104
rect 10503 7040 10519 7104
rect 10583 7040 10599 7104
rect 10663 7040 10679 7104
rect 10743 7040 10751 7104
rect 10431 6016 10751 7040
rect 10431 5952 10439 6016
rect 10503 5952 10519 6016
rect 10583 5952 10599 6016
rect 10663 5952 10679 6016
rect 10743 5952 10751 6016
rect 10431 4928 10751 5952
rect 10431 4864 10439 4928
rect 10503 4864 10519 4928
rect 10583 4864 10599 4928
rect 10663 4864 10679 4928
rect 10743 4864 10751 4928
rect 10431 4130 10751 4864
rect 10431 3894 10473 4130
rect 10709 3894 10751 4130
rect 10431 3840 10751 3894
rect 10431 3776 10439 3840
rect 10503 3776 10519 3840
rect 10583 3776 10599 3840
rect 10663 3776 10679 3840
rect 10743 3776 10751 3840
rect 10431 2752 10751 3776
rect 10431 2688 10439 2752
rect 10503 2688 10519 2752
rect 10583 2688 10599 2752
rect 10663 2688 10679 2752
rect 10743 2688 10751 2752
rect 10431 2128 10751 2688
rect 11091 16352 11411 16912
rect 11091 16288 11099 16352
rect 11163 16288 11179 16352
rect 11243 16288 11259 16352
rect 11323 16288 11339 16352
rect 11403 16288 11411 16352
rect 11091 15806 11411 16288
rect 11091 15570 11133 15806
rect 11369 15570 11411 15806
rect 11091 15264 11411 15570
rect 11091 15200 11099 15264
rect 11163 15200 11179 15264
rect 11243 15200 11259 15264
rect 11323 15200 11339 15264
rect 11403 15200 11411 15264
rect 11091 14176 11411 15200
rect 11091 14112 11099 14176
rect 11163 14112 11179 14176
rect 11243 14112 11259 14176
rect 11323 14112 11339 14176
rect 11403 14112 11411 14176
rect 11091 13088 11411 14112
rect 11091 13024 11099 13088
rect 11163 13024 11179 13088
rect 11243 13024 11259 13088
rect 11323 13024 11339 13088
rect 11403 13024 11411 13088
rect 11091 12134 11411 13024
rect 11091 12000 11133 12134
rect 11369 12000 11411 12134
rect 11091 11936 11099 12000
rect 11403 11936 11411 12000
rect 11091 11898 11133 11936
rect 11369 11898 11411 11936
rect 11091 10912 11411 11898
rect 14226 16896 14546 16912
rect 14226 16832 14234 16896
rect 14298 16832 14314 16896
rect 14378 16832 14394 16896
rect 14458 16832 14474 16896
rect 14538 16832 14546 16896
rect 14226 15808 14546 16832
rect 14226 15744 14234 15808
rect 14298 15744 14314 15808
rect 14378 15744 14394 15808
rect 14458 15744 14474 15808
rect 14538 15744 14546 15808
rect 14226 15146 14546 15744
rect 14226 14910 14268 15146
rect 14504 14910 14546 15146
rect 14226 14720 14546 14910
rect 14226 14656 14234 14720
rect 14298 14656 14314 14720
rect 14378 14656 14394 14720
rect 14458 14656 14474 14720
rect 14538 14656 14546 14720
rect 14226 13632 14546 14656
rect 14226 13568 14234 13632
rect 14298 13568 14314 13632
rect 14378 13568 14394 13632
rect 14458 13568 14474 13632
rect 14538 13568 14546 13632
rect 14226 12544 14546 13568
rect 14226 12480 14234 12544
rect 14298 12480 14314 12544
rect 14378 12480 14394 12544
rect 14458 12480 14474 12544
rect 14538 12480 14546 12544
rect 13675 11660 13741 11661
rect 13675 11596 13676 11660
rect 13740 11596 13741 11660
rect 13675 11595 13741 11596
rect 11091 10848 11099 10912
rect 11163 10848 11179 10912
rect 11243 10848 11259 10912
rect 11323 10848 11339 10912
rect 11403 10848 11411 10912
rect 11091 9824 11411 10848
rect 11091 9760 11099 9824
rect 11163 9760 11179 9824
rect 11243 9760 11259 9824
rect 11323 9760 11339 9824
rect 11403 9760 11411 9824
rect 11091 8736 11411 9760
rect 13678 9621 13738 11595
rect 14226 11474 14546 12480
rect 14226 11456 14268 11474
rect 14504 11456 14546 11474
rect 14226 11392 14234 11456
rect 14538 11392 14546 11456
rect 14226 11238 14268 11392
rect 14504 11238 14546 11392
rect 14226 10368 14546 11238
rect 14226 10304 14234 10368
rect 14298 10304 14314 10368
rect 14378 10304 14394 10368
rect 14458 10304 14474 10368
rect 14538 10304 14546 10368
rect 13675 9620 13741 9621
rect 13675 9556 13676 9620
rect 13740 9556 13741 9620
rect 13675 9555 13741 9556
rect 11091 8672 11099 8736
rect 11163 8672 11179 8736
rect 11243 8672 11259 8736
rect 11323 8672 11339 8736
rect 11403 8672 11411 8736
rect 11091 8462 11411 8672
rect 11091 8226 11133 8462
rect 11369 8226 11411 8462
rect 11091 7648 11411 8226
rect 11091 7584 11099 7648
rect 11163 7584 11179 7648
rect 11243 7584 11259 7648
rect 11323 7584 11339 7648
rect 11403 7584 11411 7648
rect 11091 6560 11411 7584
rect 11091 6496 11099 6560
rect 11163 6496 11179 6560
rect 11243 6496 11259 6560
rect 11323 6496 11339 6560
rect 11403 6496 11411 6560
rect 11091 5472 11411 6496
rect 11091 5408 11099 5472
rect 11163 5408 11179 5472
rect 11243 5408 11259 5472
rect 11323 5408 11339 5472
rect 11403 5408 11411 5472
rect 11091 4790 11411 5408
rect 11091 4554 11133 4790
rect 11369 4554 11411 4790
rect 11091 4384 11411 4554
rect 11091 4320 11099 4384
rect 11163 4320 11179 4384
rect 11243 4320 11259 4384
rect 11323 4320 11339 4384
rect 11403 4320 11411 4384
rect 11091 3296 11411 4320
rect 11091 3232 11099 3296
rect 11163 3232 11179 3296
rect 11243 3232 11259 3296
rect 11323 3232 11339 3296
rect 11403 3232 11411 3296
rect 11091 2208 11411 3232
rect 11091 2144 11099 2208
rect 11163 2144 11179 2208
rect 11243 2144 11259 2208
rect 11323 2144 11339 2208
rect 11403 2144 11411 2208
rect 11091 2128 11411 2144
rect 14226 9280 14546 10304
rect 14226 9216 14234 9280
rect 14298 9216 14314 9280
rect 14378 9216 14394 9280
rect 14458 9216 14474 9280
rect 14538 9216 14546 9280
rect 14226 8192 14546 9216
rect 14226 8128 14234 8192
rect 14298 8128 14314 8192
rect 14378 8128 14394 8192
rect 14458 8128 14474 8192
rect 14538 8128 14546 8192
rect 14226 7802 14546 8128
rect 14226 7566 14268 7802
rect 14504 7566 14546 7802
rect 14226 7104 14546 7566
rect 14226 7040 14234 7104
rect 14298 7040 14314 7104
rect 14378 7040 14394 7104
rect 14458 7040 14474 7104
rect 14538 7040 14546 7104
rect 14226 6016 14546 7040
rect 14226 5952 14234 6016
rect 14298 5952 14314 6016
rect 14378 5952 14394 6016
rect 14458 5952 14474 6016
rect 14538 5952 14546 6016
rect 14226 4928 14546 5952
rect 14226 4864 14234 4928
rect 14298 4864 14314 4928
rect 14378 4864 14394 4928
rect 14458 4864 14474 4928
rect 14538 4864 14546 4928
rect 14226 4130 14546 4864
rect 14226 3894 14268 4130
rect 14504 3894 14546 4130
rect 14226 3840 14546 3894
rect 14226 3776 14234 3840
rect 14298 3776 14314 3840
rect 14378 3776 14394 3840
rect 14458 3776 14474 3840
rect 14538 3776 14546 3840
rect 14226 2752 14546 3776
rect 14226 2688 14234 2752
rect 14298 2688 14314 2752
rect 14378 2688 14394 2752
rect 14458 2688 14474 2752
rect 14538 2688 14546 2752
rect 14226 2128 14546 2688
rect 14886 16352 15206 16912
rect 14886 16288 14894 16352
rect 14958 16288 14974 16352
rect 15038 16288 15054 16352
rect 15118 16288 15134 16352
rect 15198 16288 15206 16352
rect 14886 15806 15206 16288
rect 14886 15570 14928 15806
rect 15164 15570 15206 15806
rect 14886 15264 15206 15570
rect 14886 15200 14894 15264
rect 14958 15200 14974 15264
rect 15038 15200 15054 15264
rect 15118 15200 15134 15264
rect 15198 15200 15206 15264
rect 14886 14176 15206 15200
rect 14886 14112 14894 14176
rect 14958 14112 14974 14176
rect 15038 14112 15054 14176
rect 15118 14112 15134 14176
rect 15198 14112 15206 14176
rect 14886 13088 15206 14112
rect 14886 13024 14894 13088
rect 14958 13024 14974 13088
rect 15038 13024 15054 13088
rect 15118 13024 15134 13088
rect 15198 13024 15206 13088
rect 14886 12134 15206 13024
rect 14886 12000 14928 12134
rect 15164 12000 15206 12134
rect 14886 11936 14894 12000
rect 15198 11936 15206 12000
rect 14886 11898 14928 11936
rect 15164 11898 15206 11936
rect 14886 10912 15206 11898
rect 14886 10848 14894 10912
rect 14958 10848 14974 10912
rect 15038 10848 15054 10912
rect 15118 10848 15134 10912
rect 15198 10848 15206 10912
rect 14886 9824 15206 10848
rect 14886 9760 14894 9824
rect 14958 9760 14974 9824
rect 15038 9760 15054 9824
rect 15118 9760 15134 9824
rect 15198 9760 15206 9824
rect 14886 8736 15206 9760
rect 14886 8672 14894 8736
rect 14958 8672 14974 8736
rect 15038 8672 15054 8736
rect 15118 8672 15134 8736
rect 15198 8672 15206 8736
rect 14886 8462 15206 8672
rect 14886 8226 14928 8462
rect 15164 8226 15206 8462
rect 14886 7648 15206 8226
rect 14886 7584 14894 7648
rect 14958 7584 14974 7648
rect 15038 7584 15054 7648
rect 15118 7584 15134 7648
rect 15198 7584 15206 7648
rect 14886 6560 15206 7584
rect 14886 6496 14894 6560
rect 14958 6496 14974 6560
rect 15038 6496 15054 6560
rect 15118 6496 15134 6560
rect 15198 6496 15206 6560
rect 14886 5472 15206 6496
rect 14886 5408 14894 5472
rect 14958 5408 14974 5472
rect 15038 5408 15054 5472
rect 15118 5408 15134 5472
rect 15198 5408 15206 5472
rect 14886 4790 15206 5408
rect 14886 4554 14928 4790
rect 15164 4554 15206 4790
rect 14886 4384 15206 4554
rect 14886 4320 14894 4384
rect 14958 4320 14974 4384
rect 15038 4320 15054 4384
rect 15118 4320 15134 4384
rect 15198 4320 15206 4384
rect 14886 3296 15206 4320
rect 14886 3232 14894 3296
rect 14958 3232 14974 3296
rect 15038 3232 15054 3296
rect 15118 3232 15134 3296
rect 15198 3232 15206 3296
rect 14886 2208 15206 3232
rect 14886 2144 14894 2208
rect 14958 2144 14974 2208
rect 15038 2144 15054 2208
rect 15118 2144 15134 2208
rect 15198 2144 15206 2208
rect 14886 2128 15206 2144
<< via4 >>
rect 2883 14910 3119 15146
rect 2883 11456 3119 11474
rect 2883 11392 2913 11456
rect 2913 11392 2929 11456
rect 2929 11392 2993 11456
rect 2993 11392 3009 11456
rect 3009 11392 3073 11456
rect 3073 11392 3089 11456
rect 3089 11392 3119 11456
rect 2883 11238 3119 11392
rect 2883 7566 3119 7802
rect 2883 3894 3119 4130
rect 3543 15570 3779 15806
rect 3543 12000 3779 12134
rect 3543 11936 3573 12000
rect 3573 11936 3589 12000
rect 3589 11936 3653 12000
rect 3653 11936 3669 12000
rect 3669 11936 3733 12000
rect 3733 11936 3749 12000
rect 3749 11936 3779 12000
rect 3543 11898 3779 11936
rect 3543 8226 3779 8462
rect 3543 4554 3779 4790
rect 6678 14910 6914 15146
rect 6678 11456 6914 11474
rect 6678 11392 6708 11456
rect 6708 11392 6724 11456
rect 6724 11392 6788 11456
rect 6788 11392 6804 11456
rect 6804 11392 6868 11456
rect 6868 11392 6884 11456
rect 6884 11392 6914 11456
rect 6678 11238 6914 11392
rect 6678 7566 6914 7802
rect 6678 3894 6914 4130
rect 7338 15570 7574 15806
rect 7338 12000 7574 12134
rect 7338 11936 7368 12000
rect 7368 11936 7384 12000
rect 7384 11936 7448 12000
rect 7448 11936 7464 12000
rect 7464 11936 7528 12000
rect 7528 11936 7544 12000
rect 7544 11936 7574 12000
rect 7338 11898 7574 11936
rect 7338 8226 7574 8462
rect 7338 4554 7574 4790
rect 10473 14910 10709 15146
rect 10473 11456 10709 11474
rect 10473 11392 10503 11456
rect 10503 11392 10519 11456
rect 10519 11392 10583 11456
rect 10583 11392 10599 11456
rect 10599 11392 10663 11456
rect 10663 11392 10679 11456
rect 10679 11392 10709 11456
rect 10473 11238 10709 11392
rect 10473 7566 10709 7802
rect 10473 3894 10709 4130
rect 11133 15570 11369 15806
rect 11133 12000 11369 12134
rect 11133 11936 11163 12000
rect 11163 11936 11179 12000
rect 11179 11936 11243 12000
rect 11243 11936 11259 12000
rect 11259 11936 11323 12000
rect 11323 11936 11339 12000
rect 11339 11936 11369 12000
rect 11133 11898 11369 11936
rect 14268 14910 14504 15146
rect 14268 11456 14504 11474
rect 14268 11392 14298 11456
rect 14298 11392 14314 11456
rect 14314 11392 14378 11456
rect 14378 11392 14394 11456
rect 14394 11392 14458 11456
rect 14458 11392 14474 11456
rect 14474 11392 14504 11456
rect 14268 11238 14504 11392
rect 11133 8226 11369 8462
rect 11133 4554 11369 4790
rect 14268 7566 14504 7802
rect 14268 3894 14504 4130
rect 14928 15570 15164 15806
rect 14928 12000 15164 12134
rect 14928 11936 14958 12000
rect 14958 11936 14974 12000
rect 14974 11936 15038 12000
rect 15038 11936 15054 12000
rect 15054 11936 15118 12000
rect 15118 11936 15134 12000
rect 15134 11936 15164 12000
rect 14928 11898 15164 11936
rect 14928 8226 15164 8462
rect 14928 4554 15164 4790
<< metal5 >>
rect 1056 15806 16332 15848
rect 1056 15570 3543 15806
rect 3779 15570 7338 15806
rect 7574 15570 11133 15806
rect 11369 15570 14928 15806
rect 15164 15570 16332 15806
rect 1056 15528 16332 15570
rect 1056 15146 16332 15188
rect 1056 14910 2883 15146
rect 3119 14910 6678 15146
rect 6914 14910 10473 15146
rect 10709 14910 14268 15146
rect 14504 14910 16332 15146
rect 1056 14868 16332 14910
rect 1056 12134 16332 12176
rect 1056 11898 3543 12134
rect 3779 11898 7338 12134
rect 7574 11898 11133 12134
rect 11369 11898 14928 12134
rect 15164 11898 16332 12134
rect 1056 11856 16332 11898
rect 1056 11474 16332 11516
rect 1056 11238 2883 11474
rect 3119 11238 6678 11474
rect 6914 11238 10473 11474
rect 10709 11238 14268 11474
rect 14504 11238 16332 11474
rect 1056 11196 16332 11238
rect 1056 8462 16332 8504
rect 1056 8226 3543 8462
rect 3779 8226 7338 8462
rect 7574 8226 11133 8462
rect 11369 8226 14928 8462
rect 15164 8226 16332 8462
rect 1056 8184 16332 8226
rect 1056 7802 16332 7844
rect 1056 7566 2883 7802
rect 3119 7566 6678 7802
rect 6914 7566 10473 7802
rect 10709 7566 14268 7802
rect 14504 7566 16332 7802
rect 1056 7524 16332 7566
rect 1056 4790 16332 4832
rect 1056 4554 3543 4790
rect 3779 4554 7338 4790
rect 7574 4554 11133 4790
rect 11369 4554 14928 4790
rect 15164 4554 16332 4790
rect 1056 4512 16332 4554
rect 1056 4130 16332 4172
rect 1056 3894 2883 4130
rect 3119 3894 6678 4130
rect 6914 3894 10473 4130
rect 10709 3894 14268 4130
rect 14504 3894 16332 4130
rect 1056 3852 16332 3894
use sky130_fd_sc_hd__clkbuf_4  _120_
timestamp 0
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 0
transform -1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _122_
timestamp 0
transform -1 0 10580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _123_
timestamp 0
transform -1 0 12880 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _124_
timestamp 0
transform -1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _125_
timestamp 0
transform -1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 0
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 0
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _128_
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _129_
timestamp 0
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _130_
timestamp 0
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _131_
timestamp 0
transform -1 0 4324 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 0
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _133_
timestamp 0
transform -1 0 2944 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _134_
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _135_
timestamp 0
transform -1 0 7544 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _136_
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _138_
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _141_
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _142_
timestamp 0
transform -1 0 8740 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 0
transform -1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _144_
timestamp 0
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 0
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 0
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _148_
timestamp 0
transform -1 0 9384 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _149_
timestamp 0
transform 1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 0
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _151_
timestamp 0
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _152_
timestamp 0
transform -1 0 8832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _154_
timestamp 0
transform -1 0 2208 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp 0
transform -1 0 3312 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 0
transform 1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _157_
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 0
transform 1 0 9200 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 0
transform 1 0 9476 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 0
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 0
transform -1 0 11132 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 0
transform 1 0 10764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 0
transform -1 0 11960 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 0
transform -1 0 11408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 0
transform 1 0 13340 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 0
transform -1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 0
transform -1 0 13248 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 0
transform -1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 0
transform 1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 0
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 0
transform 1 0 11040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _174_
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _175_
timestamp 0
transform 1 0 10580 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _176_
timestamp 0
transform 1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _177_
timestamp 0
transform -1 0 2852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _178_
timestamp 0
transform 1 0 6624 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _179_
timestamp 0
transform -1 0 10120 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 0
transform -1 0 9568 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 0
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _182_
timestamp 0
transform 1 0 6624 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 0
transform 1 0 6900 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 0
transform 1 0 6440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _185_
timestamp 0
transform 1 0 9016 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 0
transform -1 0 10396 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _188_
timestamp 0
transform -1 0 8096 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp 0
transform 1 0 6808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 0
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _191_
timestamp 0
transform 1 0 6532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 0
transform 1 0 5336 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 0
transform -1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 0
transform -1 0 5244 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 0
transform 1 0 3864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _197_
timestamp 0
transform -1 0 4600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 0
transform 1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 0
transform 1 0 4324 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 0
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 0
transform 1 0 4416 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 0
transform 1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 0
transform -1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _205_
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _206_
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _207_
timestamp 0
transform -1 0 5152 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _208_
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _209_
timestamp 0
transform -1 0 11040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 0
transform -1 0 10396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 0
transform -1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _212_
timestamp 0
transform 1 0 7360 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 0
transform -1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _215_
timestamp 0
transform 1 0 11040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 0
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 0
transform 1 0 13064 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 0
transform -1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 0
transform 1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 0
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 0
transform 1 0 14260 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 0
transform -1 0 13064 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 0
transform 1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 0
transform -1 0 13432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 0
transform -1 0 14996 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 0
transform -1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 0
transform -1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 0
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 0
transform 1 0 14628 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 0
transform -1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 0
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 0
transform -1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _233_
timestamp 0
transform -1 0 11224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _234_
timestamp 0
transform 1 0 10120 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _235_
timestamp 0
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _236_
timestamp 0
transform -1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _237_
timestamp 0
transform 1 0 9200 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _238_
timestamp 0
transform 1 0 8648 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _239_
timestamp 0
transform -1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 0
transform 1 0 2024 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 0
transform 1 0 1840 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 0
transform 1 0 2024 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 0
transform 1 0 5796 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _248_
timestamp 0
transform 1 0 5428 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _249_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _250_
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 0
transform 1 0 10948 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _252_
timestamp 0
transform 1 0 8280 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _253_
timestamp 0
transform -1 0 3312 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _254_
timestamp 0
transform 1 0 7728 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _256_
timestamp 0
transform 1 0 9568 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _257_
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _258_
timestamp 0
transform 1 0 11776 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _259_
timestamp 0
transform -1 0 13984 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _260_
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _261_
timestamp 0
transform 1 0 10488 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _262_
timestamp 0
transform 1 0 2208 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 0
transform -1 0 11040 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _264_
timestamp 0
transform 1 0 5796 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _265_
timestamp 0
transform 1 0 9476 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 0
transform 1 0 6164 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _267_
timestamp 0
transform 1 0 5796 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _268_
timestamp 0
transform -1 0 6256 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 0
transform 1 0 2576 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 0
transform 1 0 1840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 0
transform 1 0 4048 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 0
transform 1 0 5796 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 0
transform -1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 0
transform -1 0 11408 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _276_
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 0
transform 1 0 12880 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 0
transform 1 0 13524 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 0
transform 1 0 13432 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 0
transform -1 0 14628 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 0
transform 1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 0
transform -1 0 3680 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 0
transform 1 0 9108 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 0
transform 1 0 9200 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _288_
timestamp 0
transform 1 0 9200 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _289_
timestamp 0
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _290_
timestamp 0
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _291_
timestamp 0
transform -1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _293_
timestamp 0
transform 1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 0
transform -1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _295_
timestamp 0
transform -1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _296_
timestamp 0
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _297_
timestamp 0
transform 1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _298_
timestamp 0
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _299_
timestamp 0
transform -1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _300_
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _301_
timestamp 0
transform -1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _302_
timestamp 0
transform -1 0 8740 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_scan_clk
timestamp 0
transform -1 0 10580 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_scan_clk
timestamp 0
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_scan_clk
timestamp 0
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_scan_clk
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_scan_clk
timestamp 0
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout5
timestamp 0
transform -1 0 3496 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout6
timestamp 0
transform 1 0 4048 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 0
transform -1 0 11132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 0
transform -1 0 10672 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18
timestamp 0
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 0
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_151
timestamp 0
transform 1 0 14996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_159
timestamp 0
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_77
timestamp 0
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_89
timestamp 0
transform 1 0 9292 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 0
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_119
timestamp 0
transform 1 0 12052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_131
timestamp 0
transform 1 0 13156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_143
timestamp 0
transform 1 0 14260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_155
timestamp 0
transform 1 0 15364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_33
timestamp 0
transform 1 0 4140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_71
timestamp 0
transform 1 0 7636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 0
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_124
timestamp 0
transform 1 0 12512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_129
timestamp 0
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_136
timestamp 0
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_161
timestamp 0
transform 1 0 15916 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_47
timestamp 0
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_67
timestamp 0
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 0
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_138
timestamp 0
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 0
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_9
timestamp 0
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_74
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_80
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_127
timestamp 0
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_161
timestamp 0
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_22
timestamp 0
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_34
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_60
timestamp 0
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_70
timestamp 0
transform 1 0 7544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_82
timestamp 0
transform 1 0 8648 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_102
timestamp 0
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_128
timestamp 0
transform 1 0 12880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_140
timestamp 0
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_152
timestamp 0
transform 1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_160
timestamp 0
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_51
timestamp 0
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_59
timestamp 0
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_67
timestamp 0
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_25
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_33
timestamp 0
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_89
timestamp 0
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_98
timestamp 0
transform 1 0 10120 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_104
timestamp 0
transform 1 0 10672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 0
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_59
timestamp 0
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_71
timestamp 0
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 0
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_113
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_125
timestamp 0
transform 1 0 12604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 0
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_161
timestamp 0
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 0
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_64
timestamp 0
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_82
timestamp 0
transform 1 0 8648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 0
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_159
timestamp 0
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_11
timestamp 0
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_33
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 0
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_107
timestamp 0
transform 1 0 10948 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_115
timestamp 0
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 0
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_161
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_78
timestamp 0
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 0
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_116
timestamp 0
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_138
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_159
timestamp 0
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 0
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_37
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_45
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 0
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_113
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_126
timestamp 0
transform 1 0 12696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 0
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_158
timestamp 0
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_49
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_66
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_76
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_44
timestamp 0
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_74
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_161
timestamp 0
transform 1 0 15916 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_11
timestamp 0
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_38
timestamp 0
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_50
timestamp 0
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_133
timestamp 0
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_155
timestamp 0
transform 1 0 15364 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_24
timestamp 0
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_49
timestamp 0
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_71
timestamp 0
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_88
timestamp 0
transform 1 0 9200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_101
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_122
timestamp 0
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_126
timestamp 0
transform 1 0 12696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_161
timestamp 0
transform 1 0 15916 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_24
timestamp 0
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_36
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_61
timestamp 0
transform 1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_72
timestamp 0
transform 1 0 7728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_104
timestamp 0
transform 1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_157
timestamp 0
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 0
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 0
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 0
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_45
timestamp 0
transform 1 0 5244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 0
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_96
timestamp 0
transform 1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_152
timestamp 0
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_31
timestamp 0
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 0
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_66
timestamp 0
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_78
timestamp 0
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_90
timestamp 0
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_102
timestamp 0
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_141
timestamp 0
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_153
timestamp 0
transform 1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 0
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_35
timestamp 0
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 0
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_113
timestamp 0
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 0
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 0
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_68
timestamp 0
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_80
timestamp 0
transform 1 0 8464 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_97
timestamp 0
transform 1 0 10028 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_103
timestamp 0
transform 1 0 10580 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_121
timestamp 0
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_143
timestamp 0
transform 1 0 14260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_155
timestamp 0
transform 1 0 15364 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_45
timestamp 0
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 0
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_108
timestamp 0
transform 1 0 11040 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_118
timestamp 0
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_161
timestamp 0
transform 1 0 15916 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_71
timestamp 0
transform 1 0 7636 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_150
timestamp 0
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 0
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 0
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_46
timestamp 0
transform 1 0 5336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_112
timestamp 0
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 0
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_149
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_161
timestamp 0
transform 1 0 15916 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_47
timestamp 0
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_60
timestamp 0
transform 1 0 6624 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_85
timestamp 0
transform 1 0 8924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_102
timestamp 0
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 0
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_121
timestamp 0
transform 1 0 12236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_133
timestamp 0
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_145
timestamp 0
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_157
timestamp 0
transform 1 0 15548 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_57
timestamp 0
transform 1 0 6348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp 0
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 0
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_93
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_98
timestamp 0
transform 1 0 10120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_110
timestamp 0
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_113
timestamp 0
transform 1 0 11500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_125
timestamp 0
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 0
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_161
timestamp 0
transform 1 0 15916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 3588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 4968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 3404 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 11776 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 9108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform 1 0 9752 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 9752 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 11224 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform 1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 15640 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 13984 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 13708 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 14904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 5888 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 0
transform -1 0 8372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 0
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 0
transform -1 0 13616 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 0
transform -1 0 14076 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 0
transform -1 0 11408 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 0
transform -1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 0
transform -1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 0
transform -1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 0
transform -1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 0
transform -1 0 14812 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 0
transform -1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 0
transform -1 0 7452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 0
transform -1 0 6716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 0
transform -1 0 11408 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 0
transform 1 0 4600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 0
transform -1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 0
transform -1 0 8372 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 0
transform -1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 0
transform -1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 0
transform -1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 0
transform -1 0 15916 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 0
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 0
transform 1 0 8832 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 0
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 0
transform -1 0 4600 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 0
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 0
transform -1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 16284 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 6256 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 11408 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
<< labels >>
rlabel metal1 s 8694 16320 8694 16320 4 VGND
rlabel metal1 s 8694 16864 8694 16864 4 VPWR
rlabel metal1 s 8326 9962 8326 9962 4 GTC.capture_en
rlabel metal1 s 1978 4148 1978 4148 4 GTC.cluster_sel\[0\]
rlabel metal1 s 4048 3978 4048 3978 4 GTC.cluster_sel\[1\]
rlabel metal1 s 7268 4794 7268 4794 4 GTC.col_addr\[0\]
rlabel metal2 s 8142 4284 8142 4284 4 GTC.col_addr\[1\]
rlabel metal2 s 6762 5440 6762 5440 4 GTC.col_addr\[2\]
rlabel metal1 s 6578 6222 6578 6222 4 GTC.col_addr\[3\]
rlabel metal1 s 2162 10200 2162 10200 4 GTC.misr_t1
rlabel metal1 s 3128 9690 3128 9690 4 GTC.misr_t2
rlabel metal1 s 2254 10030 2254 10030 4 GTC.misr_t3
rlabel metal2 s 9706 8959 9706 8959 4 GTC.mode_sel\[0\]
rlabel metal1 s 8786 10676 8786 10676 4 GTC.mode_sel\[1\]
rlabel metal1 s 3542 6630 3542 6630 4 GTC.shift_en
rlabel metal2 s 12650 4556 12650 4556 4 GTC.tier_sel\[0\]
rlabel metal1 s 11316 3570 11316 3570 4 GTC.tier_sel\[1\]
rlabel metal1 s 8924 4590 8924 4590 4 GTC.tier_sel\[2\]
rlabel metal1 s 9890 11526 9890 11526 4 TIER1.LC.scan_out
rlabel metal1 s 9660 15130 9660 15130 4 TIER1.MSS.scan_chain\[0\]
rlabel metal1 s 10534 14518 10534 14518 4 TIER1.MSS.scan_chain\[1\]
rlabel metal1 s 11500 15130 11500 15130 4 TIER1.MSS.scan_chain\[2\]
rlabel metal1 s 11454 14416 11454 14416 4 TIER1.MSS.scan_chain\[3\]
rlabel metal1 s 14398 14994 14398 14994 4 TIER1.MSS.scan_chain\[4\]
rlabel metal2 s 12190 14144 12190 14144 4 TIER1.MSS.scan_chain\[5\]
rlabel metal1 s 12880 12954 12880 12954 4 TIER1.MSS.scan_chain\[6\]
rlabel metal1 s 12052 11186 12052 11186 4 TIER1.MSS.scan_chain\[7\]
rlabel metal2 s 10902 8806 10902 8806 4 TIER1.PRAS.scan_out
rlabel metal1 s 13409 4114 13409 4114 4 TIER1.tier_sel\[0\]
rlabel metal1 s 12696 3502 12696 3502 4 TIER1.tier_sel\[1\]
rlabel metal1 s 7912 11322 7912 11322 4 TIER2.LC.scan_out
rlabel metal1 s 8142 14586 8142 14586 4 TIER2.MSS.scan_chain\[0\]
rlabel metal1 s 7498 15674 7498 15674 4 TIER2.MSS.scan_chain\[1\]
rlabel metal1 s 4876 15130 4876 15130 4 TIER2.MSS.scan_chain\[2\]
rlabel metal2 s 4370 15572 4370 15572 4 TIER2.MSS.scan_chain\[3\]
rlabel metal1 s 3956 14518 3956 14518 4 TIER2.MSS.scan_chain\[4\]
rlabel metal1 s 5750 13940 5750 13940 4 TIER2.MSS.scan_chain\[5\]
rlabel metal1 s 5842 12920 5842 12920 4 TIER2.MSS.scan_chain\[6\]
rlabel metal1 s 7222 12818 7222 12818 4 TIER2.MSS.scan_chain\[7\]
rlabel metal2 s 8510 8738 8510 8738 4 TIER2.PRAS.scan_out
rlabel metal1 s 9844 10438 9844 10438 4 TIER3.LC.scan_out
rlabel metal2 s 14674 12036 14674 12036 4 TIER3.MSS.scan_chain\[0\]
rlabel metal2 s 15870 11764 15870 11764 4 TIER3.MSS.scan_chain\[1\]
rlabel metal2 s 15318 9996 15318 9996 4 TIER3.MSS.scan_chain\[2\]
rlabel metal1 s 15226 8466 15226 8466 4 TIER3.MSS.scan_chain\[3\]
rlabel metal2 s 15870 8194 15870 8194 4 TIER3.MSS.scan_chain\[4\]
rlabel metal1 s 15870 5814 15870 5814 4 TIER3.MSS.scan_chain\[5\]
rlabel metal2 s 12834 7956 12834 7956 4 TIER3.MSS.scan_chain\[6\]
rlabel metal1 s 13524 8058 13524 8058 4 TIER3.MSS.scan_chain\[7\]
rlabel metal2 s 9982 7956 9982 7956 4 TIER3.PRAS.scan_out
rlabel metal2 s 12834 4522 12834 4522 4 _000_
rlabel metal2 s 12098 5372 12098 5372 4 _001_
rlabel metal1 s 2392 7446 2392 7446 4 _002_
rlabel metal1 s 2060 6970 2060 6970 4 _003_
rlabel metal1 s 2024 3434 2024 3434 4 _004_
rlabel metal2 s 2346 4318 2346 4318 4 _005_
rlabel metal1 s 5934 3570 5934 3570 4 _006_
rlabel metal1 s 6670 3128 6670 3128 4 _007_
rlabel metal1 s 5612 4658 5612 4658 4 _008_
rlabel metal1 s 4968 5882 4968 5882 4 _009_
rlabel metal1 s 5796 9010 5796 9010 4 _010_
rlabel metal1 s 6578 8398 6578 8398 4 _011_
rlabel metal1 s 8786 11322 8786 11322 4 _012_
rlabel metal2 s 2990 11866 2990 11866 4 _013_
rlabel metal1 s 8050 15096 8050 15096 4 _014_
rlabel metal2 s 9246 14824 9246 14824 4 _015_
rlabel metal1 s 10350 14586 10350 14586 4 _016_
rlabel metal1 s 11730 14926 11730 14926 4 _017_
rlabel metal1 s 11960 13498 11960 13498 4 _018_
rlabel metal1 s 13846 14042 13846 14042 4 _019_
rlabel metal1 s 11868 12886 11868 12886 4 _020_
rlabel metal1 s 10849 11322 10849 11322 4 _021_
rlabel metal1 s 2392 10234 2392 10234 4 _022_
rlabel metal2 s 11270 7208 11270 7208 4 _023_
rlabel metal1 s 6295 11322 6295 11322 4 _024_
rlabel metal1 s 10667 7786 10667 7786 4 _025_
rlabel metal1 s 6532 14450 6532 14450 4 _026_
rlabel metal1 s 6157 15674 6157 15674 4 _027_
rlabel metal1 s 5934 15096 5934 15096 4 _028_
rlabel metal2 s 3910 14756 3910 14756 4 _029_
rlabel metal1 s 4186 14280 4186 14280 4 _030_
rlabel metal1 s 2944 13498 2944 13498 4 _031_
rlabel metal1 s 4324 12410 4324 12410 4 _032_
rlabel metal1 s 5934 12138 5934 12138 4 _033_
rlabel metal1 s 4232 9622 4232 9622 4 _034_
rlabel metal1 s 11270 10710 11270 10710 4 _035_
rlabel metal2 s 6946 7616 6946 7616 4 _036_
rlabel metal1 s 13202 11832 13202 11832 4 _037_
rlabel metal1 s 14483 11322 14483 11322 4 _038_
rlabel metal2 s 13846 10982 13846 10982 4 _039_
rlabel metal1 s 13662 9486 13662 9486 4 _040_
rlabel metal1 s 14260 7922 14260 7922 4 _041_
rlabel metal1 s 14943 6970 14943 6970 4 _042_
rlabel metal1 s 13754 6970 13754 6970 4 _043_
rlabel metal2 s 12282 8092 12282 8092 4 _044_
rlabel metal1 s 4968 9486 4968 9486 4 _045_
rlabel metal1 s 9430 4488 9430 4488 4 _046_
rlabel metal1 s 9430 3570 9430 3570 4 _047_
rlabel metal1 s 9660 4114 9660 4114 4 _048_
rlabel metal1 s 1794 4012 1794 4012 4 _049_
rlabel metal1 s 10166 5134 10166 5134 4 _050_
rlabel metal1 s 9522 5202 9522 5202 4 _051_
rlabel metal1 s 8878 4012 8878 4012 4 _052_
rlabel metal1 s 2668 7854 2668 7854 4 _053_
rlabel metal2 s 4186 4556 4186 4556 4 _054_
rlabel metal1 s 2668 4658 2668 4658 4 _055_
rlabel metal1 s 2254 4556 2254 4556 4 _056_
rlabel metal1 s 5934 5202 5934 5202 4 _057_
rlabel metal1 s 5842 4148 5842 4148 4 _058_
rlabel metal1 s 5980 5746 5980 5746 4 _059_
rlabel metal1 s 5750 5236 5750 5236 4 _060_
rlabel metal1 s 8142 9486 8142 9486 4 _061_
rlabel metal2 s 9338 9860 9338 9860 4 _062_
rlabel metal1 s 7038 9418 7038 9418 4 _063_
rlabel metal1 s 6256 9554 6256 9554 4 _064_
rlabel metal1 s 9890 8942 9890 8942 4 _065_
rlabel metal1 s 9108 8806 9108 8806 4 _066_
rlabel metal1 s 6210 8466 6210 8466 4 _067_
rlabel metal1 s 8648 10234 8648 10234 4 _068_
rlabel metal1 s 8970 11118 8970 11118 4 _069_
rlabel metal2 s 2714 10336 2714 10336 4 _070_
rlabel metal1 s 3312 11322 3312 11322 4 _071_
rlabel metal1 s 9798 13804 9798 13804 4 _072_
rlabel metal1 s 9154 14042 9154 14042 4 _073_
rlabel metal1 s 9568 15674 9568 15674 4 _074_
rlabel metal1 s 11040 14382 11040 14382 4 _075_
rlabel metal1 s 12006 13906 12006 13906 4 _076_
rlabel metal1 s 11638 13328 11638 13328 4 _077_
rlabel metal1 s 13708 13906 13708 13906 4 _078_
rlabel metal1 s 13248 13362 13248 13362 4 _079_
rlabel metal1 s 11408 12274 11408 12274 4 _080_
rlabel metal1 s 8556 9146 8556 9146 4 _081_
rlabel metal2 s 10626 9826 10626 9826 4 _082_
rlabel metal1 s 3082 10098 3082 10098 4 _083_
rlabel metal1 s 7774 7310 7774 7310 4 _084_
rlabel metal1 s 9246 6426 9246 6426 4 _085_
rlabel metal1 s 11316 6766 11316 6766 4 _086_
rlabel metal2 s 7222 11254 7222 11254 4 _087_
rlabel metal1 s 6808 11730 6808 11730 4 _088_
rlabel metal1 s 9844 6834 9844 6834 4 _089_
rlabel metal1 s 11040 6630 11040 6630 4 _090_
rlabel metal2 s 4554 14994 4554 14994 4 _091_
rlabel metal1 s 6808 14994 6808 14994 4 _092_
rlabel metal1 s 6532 14042 6532 14042 4 _093_
rlabel metal1 s 5474 14586 5474 14586 4 _094_
rlabel metal1 s 5704 13362 5704 13362 4 _095_
rlabel metal1 s 4416 14382 4416 14382 4 _096_
rlabel metal1 s 3818 13294 3818 13294 4 _097_
rlabel metal1 s 4600 13158 4600 13158 4 _098_
rlabel metal1 s 6486 12954 6486 12954 4 _099_
rlabel metal1 s 7590 9690 7590 9690 4 _100_
rlabel metal1 s 6072 10098 6072 10098 4 _101_
rlabel metal2 s 10442 5066 10442 5066 4 _102_
rlabel metal1 s 10212 9146 10212 9146 4 _103_
rlabel metal1 s 10258 10234 10258 10234 4 _104_
rlabel metal1 s 8418 7276 8418 7276 4 _105_
rlabel metal1 s 7314 7378 7314 7378 4 _106_
rlabel metal1 s 11914 8942 11914 8942 4 _107_
rlabel metal1 s 15548 10098 15548 10098 4 _108_
rlabel metal1 s 12880 11322 12880 11322 4 _109_
rlabel metal2 s 14766 12036 14766 12036 4 _110_
rlabel metal1 s 14122 10234 14122 10234 4 _111_
rlabel metal1 s 13202 9588 13202 9588 4 _112_
rlabel metal1 s 15226 8262 15226 8262 4 _113_
rlabel metal1 s 15548 7378 15548 7378 4 _114_
rlabel metal1 s 13386 6698 13386 6698 4 _115_
rlabel metal1 s 13248 8602 13248 8602 4 _116_
rlabel metal2 s 10810 8738 10810 8738 4 _117_
rlabel metal1 s 10212 8602 10212 8602 4 _118_
rlabel metal2 s 5474 9265 5474 9265 4 _119_
rlabel metal1 s 10396 10030 10396 10030 4 clknet_0_scan_clk
rlabel metal2 s 2070 3842 2070 3842 4 clknet_2_0__leaf_scan_clk
rlabel metal1 s 2254 10710 2254 10710 4 clknet_2_1__leaf_scan_clk
rlabel metal1 s 14582 7242 14582 7242 4 clknet_2_2__leaf_scan_clk
rlabel metal1 s 9476 14926 9476 14926 4 clknet_2_3__leaf_scan_clk
rlabel metal3 s 0 14968 800 15088 4 fault_flag
port 3 nsew
rlabel metal1 s 3036 2618 3036 2618 4 net1
rlabel metal1 s 14858 9513 14858 9513 4 net10
rlabel metal1 s 4692 10030 4692 10030 4 net11
rlabel metal1 s 2760 10030 2760 10030 4 net12
rlabel metal1 s 3266 4590 3266 4590 4 net13
rlabel metal1 s 4922 9146 4922 9146 4 net14
rlabel metal1 s 3542 9010 3542 9010 4 net15
rlabel metal1 s 2208 6426 2208 6426 4 net16
rlabel metal1 s 5980 5678 5980 5678 4 net17
rlabel metal1 s 9154 4080 9154 4080 4 net18
rlabel metal1 s 11355 4794 11355 4794 4 net19
rlabel metal1 s 10166 16626 10166 16626 4 net2
rlabel metal2 s 5934 3910 5934 3910 4 net20
rlabel metal1 s 11408 3638 11408 3638 4 net21
rlabel metal1 s 6900 4182 6900 4182 4 net22
rlabel metal1 s 9292 7514 9292 7514 4 net23
rlabel metal1 s 8326 7514 8326 7514 4 net24
rlabel metal1 s 6716 5202 6716 5202 4 net25
rlabel metal2 s 9890 15674 9890 15674 4 net26
rlabel metal1 s 9430 15504 9430 15504 4 net27
rlabel metal1 s 10258 6698 10258 6698 4 net28
rlabel metal1 s 15640 8602 15640 8602 4 net29
rlabel metal1 s 14122 2482 14122 2482 4 net3
rlabel metal1 s 14122 8466 14122 8466 4 net30
rlabel metal3 s 11362 5253 11362 5253 4 net31
rlabel metal2 s 12742 13889 12742 13889 4 net32
rlabel metal1 s 12558 13294 12558 13294 4 net33
rlabel metal1 s 13340 14926 13340 14926 4 net34
rlabel metal1 s 5014 13906 5014 13906 4 net35
rlabel metal1 s 4508 12206 4508 12206 4 net36
rlabel metal1 s 7498 15130 7498 15130 4 net37
rlabel metal1 s 13708 8534 13708 8534 4 net38
rlabel metal2 s 12926 8704 12926 8704 4 net39
rlabel metal1 s 2024 12274 2024 12274 4 net4
rlabel metal2 s 13386 12410 13386 12410 4 net40
rlabel metal1 s 10994 11730 10994 11730 4 net41
rlabel metal2 s 4830 15130 4830 15130 4 net42
rlabel metal1 s 5060 13158 5060 13158 4 net43
rlabel metal1 s 11086 15538 11086 15538 4 net44
rlabel metal1 s 11684 14042 11684 14042 4 net45
rlabel metal1 s 15134 9894 15134 9894 4 net46
rlabel metal1 s 13846 12070 13846 12070 4 net47
rlabel metal1 s 15226 11594 15226 11594 4 net48
rlabel metal2 s 6762 13056 6762 13056 4 net49
rlabel metal2 s 3358 8160 3358 8160 4 net5
rlabel metal1 s 5888 13158 5888 13158 4 net50
rlabel metal1 s 10764 14042 10764 14042 4 net51
rlabel metal1 s 4692 15402 4692 15402 4 net52
rlabel metal2 s 6394 14994 6394 14994 4 net53
rlabel metal1 s 7268 11866 7268 11866 4 net54
rlabel metal1 s 4094 15470 4094 15470 4 net55
rlabel metal1 s 14904 7514 14904 7514 4 net56
rlabel metal1 s 8418 11220 8418 11220 4 net57
rlabel metal1 s 15456 6426 15456 6426 4 net58
rlabel metal1 s 13938 15130 13938 15130 4 net59
rlabel metal2 s 6486 9267 6486 9267 4 net6
rlabel metal1 s 9890 10132 9890 10132 4 net60
rlabel metal2 s 2714 11696 2714 11696 4 net61
rlabel metal1 s 3542 7514 3542 7514 4 net62
rlabel metal1 s 6019 15402 6019 15402 4 net7
rlabel metal1 s 15449 6766 15449 6766 4 net8
rlabel metal1 s 9798 15062 9798 15062 4 net9
rlabel metal2 s 46 1588 46 1588 4 reset_n
rlabel metal4 s 13708 10608 13708 10608 4 scan_clk
rlabel metal2 s 9706 17691 9706 17691 4 scan_in
rlabel metal2 s 14214 1027 14214 1027 4 test_enable
flabel metal5 s 1056 15528 16332 15848 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 11856 16332 12176 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8184 16332 8504 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4512 16332 4832 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 14886 2128 15206 16912 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 11091 2128 11411 16912 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7296 2128 7616 16912 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3501 2128 3821 16912 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 14868 16332 15188 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11196 16332 11516 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 7524 16332 7844 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3852 16332 4172 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 14226 2128 14546 16912 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10431 2128 10751 16912 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6636 2128 6956 16912 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2841 2128 3161 16912 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 400 15028 400 15028 0 FreeSans 600 0 0 0 fault_flag
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 reset_n
port 4 nsew
flabel metal3 s 16630 11568 17430 11688 0 FreeSans 600 0 0 0 scan_clk
port 5 nsew
flabel metal2 s 9678 18774 9734 19574 0 FreeSans 280 90 0 0 scan_in
port 6 nsew
flabel metal2 s 14186 0 14242 800 0 FreeSans 280 90 0 0 test_enable
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 17430 19574
<< end >>
